//  (c) Cologne Chip AG
//  FPGA Verilog netlist writer     Version: Version 4.2 (1 July 2024)
//  Compile Time: 2024-07-19 12:30:06
//  Program Run:  2024-08-22 16:24:05
//  Program Call: /home/tibrahimovic/0.git-repo/cc-toolchain-linux/cc-toolchain-linux/bin/p_r/p_r -i net/top_synth.v -o top -ccf /mnt/d/repos/LUTRAM_Stress_Test/3.build/../1.hw/constraints/constraints.ccf -cCP --verbose 
//  File Type:    Verilog

// Gatecount:   2419
module top (addr , clk , wdat , we ,
       rdat 
       ) ;

input  [7:0]addr;
input  clk;
input  [9:0]wdat;
input  we;

output [9:0]rdat;



wire [7:0]addr;
wire [9:0]wdat;
wire [9:0]rdat;
wire we;
wire clk;
wire na1_1;
wire na2_1;
wire na4_1;
wire na4_2;
wire na5_1;
wire na5_2;
wire na7_1;
wire na9_2;
wire na10_1;
wire na12_1;
wire na12_2;
wire na13_1;
wire na13_2;
wire na14_1;
wire na14_2;
wire na18_1;
wire na22_1;
wire na24_1;
wire na24_2;
wire na25_1;
wire na29_2;
wire na31_1;
wire na31_2;
wire na32_1;
wire na36_1;
wire na38_1;
wire na38_2;
wire na39_1;
wire na43_2;
wire na45_1;
wire na45_2;
wire na46_1;
wire na50_1;
wire na52_1;
wire na52_2;
wire na53_1;
wire na57_2;
wire na59_1;
wire na59_2;
wire na60_1;
wire na64_1;
wire na66_1;
wire na66_2;
wire na67_1;
wire na71_2;
wire na73_1;
wire na73_2;
wire na74_1;
wire na78_1;
wire na80_1;
wire na80_2;
wire na81_2;
wire na82_2;
wire na83_1;
wire na84_2;
wire na85_1;
wire na86_1;
wire na87_2;
wire na88_1;
wire na89_1;
wire na90_1;
wire na91_2;
wire na92_1;
wire na93_1;
wire na94_1;
wire na95_2;
wire na96_1;
wire na97_1;
wire na98_1;
wire na99_2;
wire na100_1;
wire na102_2;
wire na103_2;
wire na104_2;
wire na105_2;
wire na106_2;
wire na107_1;
wire na108_2;
wire na109_2;
wire na110_1;
wire na111_1;
wire na112_2;
wire na113_1;
wire na114_2;
wire na115_1;
wire na116_1;
wire na117_2;
wire na118_1;
wire na119_2;
wire na120_1;
wire na121_1;
wire na122_2;
wire na123_1;
wire na124_1;
wire na125_2;
wire na126_1;
wire na127_2;
wire na128_1;
wire na129_2;
wire na130_1;
wire na131_2;
wire na132_1;
wire na133_2;
wire na134_1;
wire na136_1;
wire na137_2;
wire na138_1;
wire na139_2;
wire na140_1;
wire na141_2;
wire na142_1;
wire na143_2;
wire na144_1;
wire na145_2;
wire na146_1;
wire na147_2;
wire na148_1;
wire na149_2;
wire na150_1;
wire na151_2;
wire na152_1;
wire na154_1;
wire na155_2;
wire na156_1;
wire na157_2;
wire na158_1;
wire na159_2;
wire na160_1;
wire na161_2;
wire na162_1;
wire na163_2;
wire na164_1;
wire na165_1;
wire na166_1;
wire na167_2;
wire na168_1;
wire na169_2;
wire na170_1;
wire na172_1;
wire na173_2;
wire na174_1;
wire na175_2;
wire na176_1;
wire na177_2;
wire na178_1;
wire na179_2;
wire na180_1;
wire na181_2;
wire na182_1;
wire na183_2;
wire na184_1;
wire na185_2;
wire na186_1;
wire na187_2;
wire na188_1;
wire na189_1;
wire na190_2;
wire na191_1;
wire na192_2;
wire na193_1;
wire na194_2;
wire na195_1;
wire na196_2;
wire na197_1;
wire na198_2;
wire na199_1;
wire na200_2;
wire na201_2;
wire na202_1;
wire na203_2;
wire na204_2;
wire na205_1;
wire na206_1;
wire na207_1;
wire na208_1;
wire na209_1;
wire na210_2;
wire na211_1;
wire na212_2;
wire na213_2;
wire na214_1;
wire na215_2;
wire na216_2;
wire na217_2;
wire na218_1;
wire na219_2;
wire na220_1;
wire na221_2;
wire na222_1;
wire na223_1;
wire na224_1;
wire na225_1;
wire na226_2;
wire na227_1;
wire na228_2;
wire na229_1;
wire na230_2;
wire na231_1;
wire na232_2;
wire na233_1;
wire na234_2;
wire na235_1;
wire na236_2;
wire na237_2;
wire na238_2;
wire na239_1;
wire na240_1;
wire na241_2;
wire na242_1;
wire na243_2;
wire na244_1;
wire na245_2;
wire na246_1;
wire na247_2;
wire na248_1;
wire na249_2;
wire na250_1;
wire na251_1;
wire na252_1;
wire na253_2;
wire na254_1;
wire na255_2;
wire na256_1;
wire na257_1;
wire na258_2;
wire na259_1;
wire na260_2;
wire na261_1;
wire na262_2;
wire na263_1;
wire na264_2;
wire na265_2;
wire na266_2;
wire na267_1;
wire na268_2;
wire na269_1;
wire na270_2;
wire na271_1;
wire na277_1;
wire na277_2;
wire na277_4;
wire na279_1;
wire na279_4;
wire na280_1;
wire na280_4;
wire na282_2;
wire na282_2_i;
wire na283_1;
wire na283_1_i;
wire na284_1;
wire na284_1_i;
wire na285_1;
wire na285_1_i;
wire na286_2;
wire na286_2_i;
wire na287_2;
wire na287_2_i;
wire na288_2;
wire na288_2_i;
wire na289_1;
wire na289_1_i;
wire na290_1;
wire na290_1_i;
wire na291_1;
wire na291_1_i;
wire na292_2;
wire na292_2_i;
wire na293_1;
wire na293_1_i;
wire na294_2;
wire na294_2_i;
wire na295_2;
wire na295_2_i;
wire na296_2;
wire na296_2_i;
wire na297_1;
wire na297_1_i;
wire na298_1;
wire na298_1_i;
wire na299_1;
wire na299_1_i;
wire na300_2;
wire na300_2_i;
wire na301_2;
wire na301_2_i;
wire na302_2;
wire na302_2_i;
wire na303_1;
wire na303_1_i;
wire na304_2;
wire na304_2_i;
wire na305_1;
wire na305_1_i;
wire na306_1;
wire na306_1_i;
wire na307_1;
wire na307_1_i;
wire na308_2;
wire na308_2_i;
wire na309_2;
wire na309_2_i;
wire na310_2;
wire na310_2_i;
wire na311_1;
wire na311_1_i;
wire na312_1;
wire na312_1_i;
wire na313_1;
wire na313_1_i;
wire na314_2;
wire na314_2_i;
wire na315_1;
wire na315_1_i;
wire na316_2;
wire na316_2_i;
wire na317_2;
wire na317_2_i;
wire na318_2;
wire na318_2_i;
wire na319_1;
wire na319_1_i;
wire na320_1;
wire na320_1_i;
wire na321_1;
wire na321_1_i;
wire na322_2;
wire na322_2_i;
wire na323_2;
wire na323_2_i;
wire na324_2;
wire na324_2_i;
wire na325_1;
wire na325_1_i;
wire na326_2;
wire na326_2_i;
wire na327_1;
wire na327_1_i;
wire na328_1;
wire na328_1_i;
wire na329_1;
wire na329_1_i;
wire na330_2;
wire na330_2_i;
wire na331_2;
wire na331_2_i;
wire na332_2;
wire na332_2_i;
wire na333_1;
wire na333_1_i;
wire na334_1;
wire na334_1_i;
wire na335_1;
wire na335_1_i;
wire na336_2;
wire na336_2_i;
wire na337_1;
wire na337_1_i;
wire na338_2;
wire na338_2_i;
wire na339_2;
wire na339_2_i;
wire na340_2;
wire na340_2_i;
wire na341_1;
wire na341_1_i;
wire na342_1;
wire na342_1_i;
wire na343_1;
wire na343_1_i;
wire na344_2;
wire na344_2_i;
wire na345_2;
wire na345_2_i;
wire na346_2;
wire na346_2_i;
wire na347_1;
wire na347_1_i;
wire na348_2;
wire na348_2_i;
wire na349_1;
wire na349_1_i;
wire na350_1;
wire na350_1_i;
wire na351_1;
wire na351_1_i;
wire na352_2;
wire na352_2_i;
wire na353_2;
wire na353_2_i;
wire na354_2;
wire na354_2_i;
wire na355_1;
wire na355_1_i;
wire na356_1;
wire na356_1_i;
wire na357_1;
wire na357_1_i;
wire na358_2;
wire na358_2_i;
wire na359_1;
wire na359_1_i;
wire na360_2;
wire na360_2_i;
wire na361_2;
wire na361_2_i;
wire na362_2;
wire na362_2_i;
wire na363_1;
wire na363_1_i;
wire na364_1;
wire na364_1_i;
wire na365_1;
wire na365_1_i;
wire na366_2;
wire na366_2_i;
wire na367_2;
wire na367_2_i;
wire na368_2;
wire na368_2_i;
wire na369_1;
wire na369_1_i;
wire na370_2;
wire na370_2_i;
wire na371_1;
wire na371_1_i;
wire na372_1;
wire na372_1_i;
wire na373_1;
wire na373_1_i;
wire na374_2;
wire na374_2_i;
wire na375_2;
wire na375_2_i;
wire na376_2;
wire na376_2_i;
wire na377_1;
wire na377_1_i;
wire na378_1;
wire na378_1_i;
wire na379_1;
wire na379_1_i;
wire na380_2;
wire na380_2_i;
wire na381_1;
wire na381_1_i;
wire na382_2;
wire na382_2_i;
wire na383_2;
wire na383_2_i;
wire na384_2;
wire na384_2_i;
wire na385_1;
wire na385_1_i;
wire na386_1;
wire na386_1_i;
wire na387_1;
wire na387_1_i;
wire na388_2;
wire na388_2_i;
wire na389_2;
wire na389_2_i;
wire na390_2;
wire na390_2_i;
wire na391_1;
wire na391_1_i;
wire na392_2;
wire na392_2_i;
wire na393_1;
wire na393_1_i;
wire na394_1;
wire na394_1_i;
wire na395_1;
wire na395_1_i;
wire na396_2;
wire na396_2_i;
wire na397_2;
wire na397_2_i;
wire na398_2;
wire na398_2_i;
wire na399_1;
wire na399_1_i;
wire na400_1;
wire na400_1_i;
wire na401_1;
wire na401_1_i;
wire na402_2;
wire na402_2_i;
wire na403_1;
wire na403_1_i;
wire na404_2;
wire na404_2_i;
wire na405_2;
wire na405_2_i;
wire na406_2;
wire na406_2_i;
wire na407_1;
wire na407_1_i;
wire na408_1;
wire na408_1_i;
wire na409_1;
wire na409_1_i;
wire na410_2;
wire na410_2_i;
wire na411_2;
wire na411_2_i;
wire na412_2;
wire na412_2_i;
wire na413_1;
wire na413_1_i;
wire na414_2;
wire na414_2_i;
wire na415_1;
wire na415_1_i;
wire na416_1;
wire na416_1_i;
wire na417_1;
wire na417_1_i;
wire na418_2;
wire na418_2_i;
wire na419_2;
wire na419_2_i;
wire na420_2;
wire na420_2_i;
wire na421_1;
wire na421_1_i;
wire na422_1;
wire na422_1_i;
wire na423_1;
wire na423_1_i;
wire na424_2;
wire na424_2_i;
wire na425_1;
wire na425_1_i;
wire na426_2;
wire na426_2_i;
wire na427_2;
wire na427_2_i;
wire na428_2;
wire na428_2_i;
wire na429_1;
wire na429_1_i;
wire na430_1;
wire na430_1_i;
wire na431_1;
wire na431_1_i;
wire na432_2;
wire na432_2_i;
wire na433_2;
wire na433_2_i;
wire na434_2;
wire na434_2_i;
wire na435_1;
wire na435_1_i;
wire na436_2;
wire na436_2_i;
wire na437_1;
wire na437_1_i;
wire na438_1;
wire na438_1_i;
wire na439_1;
wire na439_1_i;
wire na440_2;
wire na440_2_i;
wire na441_2;
wire na441_2_i;
wire na442_2;
wire na442_2_i;
wire na443_1;
wire na443_1_i;
wire na444_1;
wire na444_1_i;
wire na445_1;
wire na445_1_i;
wire na446_2;
wire na446_2_i;
wire na447_1;
wire na447_1_i;
wire na448_2;
wire na448_2_i;
wire na449_2;
wire na449_2_i;
wire na450_2;
wire na450_2_i;
wire na451_1;
wire na451_1_i;
wire na452_1;
wire na452_1_i;
wire na453_1;
wire na453_1_i;
wire na454_2;
wire na454_2_i;
wire na455_2;
wire na455_2_i;
wire na456_2;
wire na456_2_i;
wire na457_1;
wire na457_1_i;
wire na458_2;
wire na458_2_i;
wire na459_1;
wire na459_1_i;
wire na460_1;
wire na460_1_i;
wire na461_1;
wire na461_1_i;
wire na462_2;
wire na462_2_i;
wire na463_2;
wire na463_2_i;
wire na464_2;
wire na464_2_i;
wire na465_1;
wire na465_1_i;
wire na466_1;
wire na466_1_i;
wire na467_1;
wire na467_1_i;
wire na468_2;
wire na468_2_i;
wire na469_1;
wire na469_1_i;
wire na470_2;
wire na470_2_i;
wire na471_2;
wire na471_2_i;
wire na472_2;
wire na472_2_i;
wire na473_1;
wire na473_1_i;
wire na474_1;
wire na474_1_i;
wire na475_1;
wire na475_1_i;
wire na476_2;
wire na476_2_i;
wire na477_2;
wire na477_2_i;
wire na478_2;
wire na478_2_i;
wire na479_1;
wire na479_1_i;
wire na480_2;
wire na480_2_i;
wire na481_1;
wire na481_1_i;
wire na482_1;
wire na482_1_i;
wire na483_1;
wire na483_1_i;
wire na484_2;
wire na484_2_i;
wire na485_2;
wire na485_2_i;
wire na486_2;
wire na486_2_i;
wire na487_1;
wire na487_1_i;
wire na488_1;
wire na488_1_i;
wire na489_1;
wire na489_1_i;
wire na490_2;
wire na490_2_i;
wire na491_1;
wire na491_1_i;
wire na492_2;
wire na492_2_i;
wire na493_2;
wire na493_2_i;
wire na494_2;
wire na494_2_i;
wire na495_1;
wire na495_1_i;
wire na496_1;
wire na496_1_i;
wire na497_1;
wire na497_1_i;
wire na498_2;
wire na498_2_i;
wire na499_2;
wire na499_2_i;
wire na500_2;
wire na500_2_i;
wire na501_1;
wire na501_1_i;
wire na502_2;
wire na502_2_i;
wire na503_1;
wire na503_1_i;
wire na504_1;
wire na504_1_i;
wire na505_1;
wire na505_1_i;
wire na506_2;
wire na506_2_i;
wire na507_2;
wire na507_2_i;
wire na508_2;
wire na508_2_i;
wire na509_1;
wire na509_1_i;
wire na510_1;
wire na510_1_i;
wire na511_1;
wire na511_1_i;
wire na512_2;
wire na512_2_i;
wire na513_1;
wire na513_1_i;
wire na514_2;
wire na514_2_i;
wire na515_2;
wire na515_2_i;
wire na516_2;
wire na516_2_i;
wire na517_1;
wire na517_1_i;
wire na518_1;
wire na518_1_i;
wire na519_1;
wire na519_1_i;
wire na520_2;
wire na520_2_i;
wire na521_2;
wire na521_2_i;
wire na522_2;
wire na522_2_i;
wire na523_1;
wire na523_1_i;
wire na524_2;
wire na524_2_i;
wire na525_1;
wire na525_1_i;
wire na526_1;
wire na526_1_i;
wire na527_1;
wire na527_1_i;
wire na528_2;
wire na528_2_i;
wire na529_2;
wire na529_2_i;
wire na530_2;
wire na530_2_i;
wire na531_1;
wire na531_1_i;
wire na532_1;
wire na532_1_i;
wire na533_1;
wire na533_1_i;
wire na534_2;
wire na534_2_i;
wire na535_1;
wire na535_1_i;
wire na536_2;
wire na536_2_i;
wire na537_2;
wire na537_2_i;
wire na538_2;
wire na538_2_i;
wire na539_1;
wire na539_1_i;
wire na540_1;
wire na540_1_i;
wire na541_1;
wire na541_1_i;
wire na542_2;
wire na542_2_i;
wire na543_2;
wire na543_2_i;
wire na544_2;
wire na544_2_i;
wire na545_1;
wire na545_1_i;
wire na546_2;
wire na546_2_i;
wire na547_1;
wire na547_1_i;
wire na548_1;
wire na548_1_i;
wire na549_1;
wire na549_1_i;
wire na550_2;
wire na550_2_i;
wire na551_2;
wire na551_2_i;
wire na552_2;
wire na552_2_i;
wire na553_1;
wire na553_1_i;
wire na554_1;
wire na554_1_i;
wire na555_1;
wire na555_1_i;
wire na556_2;
wire na556_2_i;
wire na557_1;
wire na557_1_i;
wire na558_2;
wire na558_2_i;
wire na559_2;
wire na559_2_i;
wire na560_2;
wire na560_2_i;
wire na561_1;
wire na561_1_i;
wire na562_1;
wire na562_1_i;
wire na563_1;
wire na563_1_i;
wire na564_2;
wire na564_2_i;
wire na565_2;
wire na565_2_i;
wire na566_2;
wire na566_2_i;
wire na567_1;
wire na567_1_i;
wire na568_2;
wire na568_2_i;
wire na569_1;
wire na569_1_i;
wire na570_1;
wire na570_1_i;
wire na571_1;
wire na571_1_i;
wire na572_2;
wire na572_2_i;
wire na573_2;
wire na573_2_i;
wire na574_2;
wire na574_2_i;
wire na575_1;
wire na575_1_i;
wire na576_1;
wire na576_1_i;
wire na577_1;
wire na577_1_i;
wire na578_2;
wire na578_2_i;
wire na579_1;
wire na579_1_i;
wire na580_2;
wire na580_2_i;
wire na581_2;
wire na581_2_i;
wire na582_2;
wire na582_2_i;
wire na583_1;
wire na583_1_i;
wire na584_1;
wire na584_1_i;
wire na585_1;
wire na585_1_i;
wire na586_2;
wire na586_2_i;
wire na587_2;
wire na587_2_i;
wire na588_2;
wire na588_2_i;
wire na589_1;
wire na589_1_i;
wire na590_2;
wire na590_2_i;
wire na591_1;
wire na591_1_i;
wire na592_1;
wire na592_1_i;
wire na593_1;
wire na593_1_i;
wire na594_2;
wire na594_2_i;
wire na595_2;
wire na595_2_i;
wire na596_2;
wire na596_2_i;
wire na597_1;
wire na597_1_i;
wire na598_1;
wire na598_1_i;
wire na599_1;
wire na599_1_i;
wire na600_2;
wire na600_2_i;
wire na601_1;
wire na601_1_i;
wire na602_2;
wire na602_2_i;
wire na603_2;
wire na603_2_i;
wire na604_2;
wire na604_2_i;
wire na605_1;
wire na605_1_i;
wire na606_1;
wire na606_1_i;
wire na607_1;
wire na607_1_i;
wire na608_2;
wire na608_2_i;
wire na609_2;
wire na609_2_i;
wire na610_2;
wire na610_2_i;
wire na611_1;
wire na611_1_i;
wire na612_2;
wire na612_2_i;
wire na613_1;
wire na613_1_i;
wire na614_1;
wire na614_1_i;
wire na615_1;
wire na615_1_i;
wire na616_2;
wire na616_2_i;
wire na617_2;
wire na617_2_i;
wire na618_2;
wire na618_2_i;
wire na619_1;
wire na619_1_i;
wire na620_1;
wire na620_1_i;
wire na621_1;
wire na621_1_i;
wire na622_2;
wire na622_2_i;
wire na623_1;
wire na623_1_i;
wire na624_2;
wire na624_2_i;
wire na625_2;
wire na625_2_i;
wire na626_2;
wire na626_2_i;
wire na627_1;
wire na627_1_i;
wire na628_1;
wire na628_1_i;
wire na629_1;
wire na629_1_i;
wire na630_2;
wire na630_2_i;
wire na631_2;
wire na631_2_i;
wire na632_2;
wire na632_2_i;
wire na633_1;
wire na633_1_i;
wire na634_2;
wire na634_2_i;
wire na635_1;
wire na635_1_i;
wire na636_1;
wire na636_1_i;
wire na637_1;
wire na637_1_i;
wire na638_2;
wire na638_2_i;
wire na639_2;
wire na639_2_i;
wire na640_2;
wire na640_2_i;
wire na641_1;
wire na641_1_i;
wire na642_1;
wire na642_1_i;
wire na643_1;
wire na643_1_i;
wire na644_2;
wire na644_2_i;
wire na645_1;
wire na645_1_i;
wire na646_2;
wire na646_2_i;
wire na647_2;
wire na647_2_i;
wire na648_2;
wire na648_2_i;
wire na649_1;
wire na649_1_i;
wire na650_1;
wire na650_1_i;
wire na651_1;
wire na651_1_i;
wire na652_2;
wire na652_2_i;
wire na653_2;
wire na653_2_i;
wire na654_2;
wire na654_2_i;
wire na655_1;
wire na655_1_i;
wire na656_2;
wire na656_2_i;
wire na657_1;
wire na657_1_i;
wire na658_1;
wire na658_1_i;
wire na659_1;
wire na659_1_i;
wire na660_2;
wire na660_2_i;
wire na661_2;
wire na661_2_i;
wire na662_2;
wire na662_2_i;
wire na663_1;
wire na663_1_i;
wire na664_1;
wire na664_1_i;
wire na665_1;
wire na665_1_i;
wire na666_2;
wire na666_2_i;
wire na667_1;
wire na667_1_i;
wire na668_2;
wire na668_2_i;
wire na669_2;
wire na669_2_i;
wire na670_2;
wire na670_2_i;
wire na671_1;
wire na671_1_i;
wire na672_1;
wire na672_1_i;
wire na673_1;
wire na673_1_i;
wire na674_2;
wire na674_2_i;
wire na675_2;
wire na675_2_i;
wire na676_2;
wire na676_2_i;
wire na677_1;
wire na677_1_i;
wire na678_2;
wire na678_2_i;
wire na679_1;
wire na679_1_i;
wire na680_1;
wire na680_1_i;
wire na681_1;
wire na681_1_i;
wire na682_2;
wire na682_2_i;
wire na683_2;
wire na683_2_i;
wire na684_2;
wire na684_2_i;
wire na685_1;
wire na685_1_i;
wire na686_1;
wire na686_1_i;
wire na687_1;
wire na687_1_i;
wire na688_2;
wire na688_2_i;
wire na689_1;
wire na689_1_i;
wire na690_2;
wire na690_2_i;
wire na691_2;
wire na691_2_i;
wire na692_2;
wire na692_2_i;
wire na693_1;
wire na693_1_i;
wire na694_1;
wire na694_1_i;
wire na695_1;
wire na695_1_i;
wire na696_2;
wire na696_2_i;
wire na697_2;
wire na697_2_i;
wire na698_2;
wire na698_2_i;
wire na699_1;
wire na699_1_i;
wire na700_2;
wire na700_2_i;
wire na701_1;
wire na701_1_i;
wire na702_1;
wire na702_1_i;
wire na703_1;
wire na703_1_i;
wire na704_2;
wire na704_2_i;
wire na705_2;
wire na705_2_i;
wire na706_2;
wire na706_2_i;
wire na707_1;
wire na707_1_i;
wire na708_1;
wire na708_1_i;
wire na709_1;
wire na709_1_i;
wire na710_2;
wire na710_2_i;
wire na711_1;
wire na711_1_i;
wire na712_2;
wire na712_2_i;
wire na713_2;
wire na713_2_i;
wire na714_2;
wire na714_2_i;
wire na715_1;
wire na715_1_i;
wire na716_1;
wire na716_1_i;
wire na717_1;
wire na717_1_i;
wire na718_2;
wire na718_2_i;
wire na719_2;
wire na719_2_i;
wire na720_2;
wire na720_2_i;
wire na721_1;
wire na721_1_i;
wire na722_2;
wire na722_2_i;
wire na723_1;
wire na723_1_i;
wire na724_1;
wire na724_1_i;
wire na725_1;
wire na725_1_i;
wire na726_2;
wire na726_2_i;
wire na727_2;
wire na727_2_i;
wire na728_2;
wire na728_2_i;
wire na729_1;
wire na729_1_i;
wire na730_1;
wire na730_1_i;
wire na731_1;
wire na731_1_i;
wire na732_2;
wire na732_2_i;
wire na733_1;
wire na733_1_i;
wire na734_2;
wire na734_2_i;
wire na735_2;
wire na735_2_i;
wire na736_2;
wire na736_2_i;
wire na737_1;
wire na737_1_i;
wire na738_1;
wire na738_1_i;
wire na739_1;
wire na739_1_i;
wire na740_2;
wire na740_2_i;
wire na741_2;
wire na741_2_i;
wire na742_2;
wire na742_2_i;
wire na743_1;
wire na743_1_i;
wire na744_2;
wire na744_2_i;
wire na745_1;
wire na745_1_i;
wire na746_1;
wire na746_1_i;
wire na747_1;
wire na747_1_i;
wire na748_2;
wire na748_2_i;
wire na749_2;
wire na749_2_i;
wire na750_2;
wire na750_2_i;
wire na751_1;
wire na751_1_i;
wire na752_1;
wire na752_1_i;
wire na753_1;
wire na753_1_i;
wire na754_2;
wire na754_2_i;
wire na755_1;
wire na755_1_i;
wire na756_2;
wire na756_2_i;
wire na757_2;
wire na757_2_i;
wire na758_2;
wire na758_2_i;
wire na759_1;
wire na759_1_i;
wire na760_1;
wire na760_1_i;
wire na761_1;
wire na761_1_i;
wire na762_2;
wire na762_2_i;
wire na763_2;
wire na763_2_i;
wire na764_2;
wire na764_2_i;
wire na765_1;
wire na765_1_i;
wire na766_2;
wire na766_2_i;
wire na767_1;
wire na767_1_i;
wire na768_1;
wire na768_1_i;
wire na769_1;
wire na769_1_i;
wire na770_2;
wire na770_2_i;
wire na771_2;
wire na771_2_i;
wire na772_2;
wire na772_2_i;
wire na773_1;
wire na773_1_i;
wire na774_1;
wire na774_1_i;
wire na775_1;
wire na775_1_i;
wire na776_2;
wire na776_2_i;
wire na777_1;
wire na777_1_i;
wire na778_2;
wire na778_2_i;
wire na779_2;
wire na779_2_i;
wire na780_2;
wire na780_2_i;
wire na781_1;
wire na781_1_i;
wire na782_1;
wire na782_1_i;
wire na783_1;
wire na783_1_i;
wire na784_2;
wire na784_2_i;
wire na785_2;
wire na785_2_i;
wire na786_2;
wire na786_2_i;
wire na787_1;
wire na787_1_i;
wire na788_2;
wire na788_2_i;
wire na789_1;
wire na789_1_i;
wire na790_1;
wire na790_1_i;
wire na791_1;
wire na791_1_i;
wire na792_2;
wire na792_2_i;
wire na793_2;
wire na793_2_i;
wire na794_2;
wire na794_2_i;
wire na795_1;
wire na795_1_i;
wire na796_1;
wire na796_1_i;
wire na797_1;
wire na797_1_i;
wire na798_2;
wire na798_2_i;
wire na799_1;
wire na799_1_i;
wire na800_2;
wire na800_2_i;
wire na801_2;
wire na801_2_i;
wire na802_2;
wire na802_2_i;
wire na803_1;
wire na803_1_i;
wire na804_1;
wire na804_1_i;
wire na805_1;
wire na805_1_i;
wire na806_2;
wire na806_2_i;
wire na807_2;
wire na807_2_i;
wire na808_2;
wire na808_2_i;
wire na809_1;
wire na809_1_i;
wire na810_2;
wire na810_2_i;
wire na811_1;
wire na811_1_i;
wire na812_1;
wire na812_1_i;
wire na813_1;
wire na813_1_i;
wire na814_2;
wire na814_2_i;
wire na815_2;
wire na815_2_i;
wire na816_2;
wire na816_2_i;
wire na817_1;
wire na817_1_i;
wire na818_1;
wire na818_1_i;
wire na819_1;
wire na819_1_i;
wire na820_2;
wire na820_2_i;
wire na821_1;
wire na821_1_i;
wire na822_2;
wire na822_2_i;
wire na823_2;
wire na823_2_i;
wire na824_2;
wire na824_2_i;
wire na825_1;
wire na825_1_i;
wire na826_1;
wire na826_1_i;
wire na827_1;
wire na827_1_i;
wire na828_2;
wire na828_2_i;
wire na829_2;
wire na829_2_i;
wire na830_2;
wire na830_2_i;
wire na831_1;
wire na831_1_i;
wire na832_2;
wire na832_2_i;
wire na833_1;
wire na833_1_i;
wire na834_1;
wire na834_1_i;
wire na835_1;
wire na835_1_i;
wire na836_2;
wire na836_2_i;
wire na837_2;
wire na837_2_i;
wire na838_2;
wire na838_2_i;
wire na839_1;
wire na839_1_i;
wire na840_1;
wire na840_1_i;
wire na841_1;
wire na841_1_i;
wire na842_2;
wire na842_2_i;
wire na843_1;
wire na843_1_i;
wire na844_2;
wire na844_2_i;
wire na845_2;
wire na845_2_i;
wire na846_2;
wire na846_2_i;
wire na847_1;
wire na847_1_i;
wire na848_1;
wire na848_1_i;
wire na849_1;
wire na849_1_i;
wire na850_2;
wire na850_2_i;
wire na851_2;
wire na851_2_i;
wire na852_2;
wire na852_2_i;
wire na853_1;
wire na853_1_i;
wire na854_2;
wire na854_2_i;
wire na855_1;
wire na855_1_i;
wire na856_1;
wire na856_1_i;
wire na857_1;
wire na857_1_i;
wire na858_2;
wire na858_2_i;
wire na859_2;
wire na859_2_i;
wire na860_2;
wire na860_2_i;
wire na861_1;
wire na861_1_i;
wire na862_1;
wire na862_1_i;
wire na863_1;
wire na863_1_i;
wire na864_2;
wire na864_2_i;
wire na865_1;
wire na865_1_i;
wire na866_2;
wire na866_2_i;
wire na867_2;
wire na867_2_i;
wire na868_2;
wire na868_2_i;
wire na869_1;
wire na869_1_i;
wire na870_1;
wire na870_1_i;
wire na871_1;
wire na871_1_i;
wire na872_2;
wire na872_2_i;
wire na873_2;
wire na873_2_i;
wire na874_2;
wire na874_2_i;
wire na875_1;
wire na875_1_i;
wire na876_2;
wire na876_2_i;
wire na877_1;
wire na877_1_i;
wire na878_1;
wire na878_1_i;
wire na879_1;
wire na879_1_i;
wire na880_2;
wire na880_2_i;
wire na881_2;
wire na881_2_i;
wire na882_2;
wire na882_2_i;
wire na883_1;
wire na883_1_i;
wire na884_1;
wire na884_1_i;
wire na885_1;
wire na885_1_i;
wire na886_2;
wire na886_2_i;
wire na887_1;
wire na887_1_i;
wire na888_2;
wire na888_2_i;
wire na889_2;
wire na889_2_i;
wire na890_2;
wire na890_2_i;
wire na891_1;
wire na891_1_i;
wire na892_1;
wire na892_1_i;
wire na893_1;
wire na893_1_i;
wire na894_2;
wire na894_2_i;
wire na895_2;
wire na895_2_i;
wire na896_2;
wire na896_2_i;
wire na897_1;
wire na897_1_i;
wire na898_2;
wire na898_2_i;
wire na899_1;
wire na899_1_i;
wire na900_1;
wire na900_1_i;
wire na901_1;
wire na901_1_i;
wire na902_2;
wire na902_2_i;
wire na903_2;
wire na903_2_i;
wire na904_2;
wire na904_2_i;
wire na905_1;
wire na905_1_i;
wire na906_1;
wire na906_1_i;
wire na907_1;
wire na907_1_i;
wire na908_2;
wire na908_2_i;
wire na909_1;
wire na909_1_i;
wire na910_2;
wire na910_2_i;
wire na911_2;
wire na911_2_i;
wire na912_2;
wire na912_2_i;
wire na913_1;
wire na913_1_i;
wire na914_1;
wire na914_1_i;
wire na915_1;
wire na915_1_i;
wire na916_2;
wire na916_2_i;
wire na917_2;
wire na917_2_i;
wire na918_2;
wire na918_2_i;
wire na919_1;
wire na919_1_i;
wire na920_2;
wire na920_2_i;
wire na921_1;
wire na921_1_i;
wire na922_1;
wire na922_1_i;
wire na923_1;
wire na923_1_i;
wire na924_2;
wire na924_2_i;
wire na925_2;
wire na925_2_i;
wire na926_2;
wire na926_2_i;
wire na927_1;
wire na927_1_i;
wire na928_1;
wire na928_1_i;
wire na929_1;
wire na929_1_i;
wire na930_2;
wire na930_2_i;
wire na931_1;
wire na931_1_i;
wire na932_2;
wire na932_2_i;
wire na933_2;
wire na933_2_i;
wire na934_2;
wire na934_2_i;
wire na935_1;
wire na935_1_i;
wire na936_1;
wire na936_1_i;
wire na937_1;
wire na937_1_i;
wire na938_2;
wire na938_2_i;
wire na939_2;
wire na939_2_i;
wire na940_2;
wire na940_2_i;
wire na941_1;
wire na941_1_i;
wire na942_2;
wire na942_2_i;
wire na943_1;
wire na943_1_i;
wire na944_1;
wire na944_1_i;
wire na945_1;
wire na945_1_i;
wire na946_2;
wire na946_2_i;
wire na947_2;
wire na947_2_i;
wire na948_2;
wire na948_2_i;
wire na949_1;
wire na949_1_i;
wire na950_1;
wire na950_1_i;
wire na951_1;
wire na951_1_i;
wire na952_2;
wire na952_2_i;
wire na953_1;
wire na953_1_i;
wire na954_2;
wire na954_2_i;
wire na955_2;
wire na955_2_i;
wire na956_2;
wire na956_2_i;
wire na957_1;
wire na957_1_i;
wire na958_1;
wire na958_1_i;
wire na959_1;
wire na959_1_i;
wire na960_2;
wire na960_2_i;
wire na961_2;
wire na961_2_i;
wire na962_2;
wire na962_2_i;
wire na963_1;
wire na963_1_i;
wire na964_2;
wire na964_2_i;
wire na965_1;
wire na965_1_i;
wire na966_1;
wire na966_1_i;
wire na967_1;
wire na967_1_i;
wire na968_2;
wire na968_2_i;
wire na969_2;
wire na969_2_i;
wire na970_2;
wire na970_2_i;
wire na971_1;
wire na971_1_i;
wire na972_1;
wire na972_1_i;
wire na973_1;
wire na973_1_i;
wire na974_2;
wire na974_2_i;
wire na975_1;
wire na975_1_i;
wire na976_2;
wire na976_2_i;
wire na977_2;
wire na977_2_i;
wire na978_2;
wire na978_2_i;
wire na979_1;
wire na979_1_i;
wire na980_1;
wire na980_1_i;
wire na981_1;
wire na981_1_i;
wire na982_2;
wire na982_2_i;
wire na983_2;
wire na983_2_i;
wire na984_2;
wire na984_2_i;
wire na985_1;
wire na985_1_i;
wire na986_1;
wire na986_1_i;
wire na987_1;
wire na987_1_i;
wire na988_2;
wire na988_2_i;
wire na989_1;
wire na989_1_i;
wire na990_2;
wire na990_2_i;
wire na991_1;
wire na991_1_i;
wire na992_2;
wire na992_2_i;
wire na993_2;
wire na993_2_i;
wire na994_2;
wire na994_2_i;
wire na995_1;
wire na995_1_i;
wire na996_2;
wire na996_2_i;
wire na997_1;
wire na997_1_i;
wire na998_2;
wire na998_2_i;
wire na999_1;
wire na999_1_i;
wire na1000_1;
wire na1000_1_i;
wire na1001_1;
wire na1001_1_i;
wire na1002_2;
wire na1002_2_i;
wire na1003_1;
wire na1003_1_i;
wire na1004_2;
wire na1004_2_i;
wire na1005_1;
wire na1005_1_i;
wire na1006_2;
wire na1006_2_i;
wire na1007_2;
wire na1007_2_i;
wire na1008_2;
wire na1008_2_i;
wire na1009_1;
wire na1009_1_i;
wire na1010_2;
wire na1010_2_i;
wire na1011_1;
wire na1011_1_i;
wire na1012_2;
wire na1012_2_i;
wire na1013_1;
wire na1013_1_i;
wire na1014_1;
wire na1014_1_i;
wire na1015_1;
wire na1015_1_i;
wire na1016_2;
wire na1016_2_i;
wire na1017_1;
wire na1017_1_i;
wire na1018_2;
wire na1018_2_i;
wire na1019_1;
wire na1019_1_i;
wire na1020_2;
wire na1020_2_i;
wire na1021_2;
wire na1021_2_i;
wire na1022_2;
wire na1022_2_i;
wire na1023_1;
wire na1023_1_i;
wire na1024_2;
wire na1024_2_i;
wire na1025_1;
wire na1025_1_i;
wire na1026_2;
wire na1026_2_i;
wire na1027_1;
wire na1027_1_i;
wire na1028_1;
wire na1028_1_i;
wire na1029_1;
wire na1029_1_i;
wire na1030_2;
wire na1030_2_i;
wire na1031_1;
wire na1031_1_i;
wire na1032_2;
wire na1032_2_i;
wire na1033_1;
wire na1033_1_i;
wire na1034_2;
wire na1034_2_i;
wire na1035_2;
wire na1035_2_i;
wire na1036_2;
wire na1036_2_i;
wire na1037_1;
wire na1037_1_i;
wire na1038_2;
wire na1038_2_i;
wire na1039_1;
wire na1039_1_i;
wire na1040_2;
wire na1040_2_i;
wire na1041_1;
wire na1041_1_i;
wire na1042_1;
wire na1042_1_i;
wire na1043_1;
wire na1043_1_i;
wire na1044_2;
wire na1044_2_i;
wire na1045_1;
wire na1045_1_i;
wire na1046_2;
wire na1046_2_i;
wire na1047_1;
wire na1047_1_i;
wire na1048_2;
wire na1048_2_i;
wire na1049_2;
wire na1049_2_i;
wire na1050_2;
wire na1050_2_i;
wire na1051_1;
wire na1051_1_i;
wire na1052_2;
wire na1052_2_i;
wire na1053_1;
wire na1053_1_i;
wire na1054_2;
wire na1054_2_i;
wire na1055_1;
wire na1055_1_i;
wire na1056_1;
wire na1056_1_i;
wire na1057_1;
wire na1057_1_i;
wire na1058_2;
wire na1058_2_i;
wire na1059_1;
wire na1059_1_i;
wire na1060_2;
wire na1060_2_i;
wire na1061_1;
wire na1061_1_i;
wire na1062_2;
wire na1062_2_i;
wire na1063_2;
wire na1063_2_i;
wire na1064_2;
wire na1064_2_i;
wire na1065_1;
wire na1065_1_i;
wire na1066_2;
wire na1066_2_i;
wire na1067_1;
wire na1067_1_i;
wire na1068_2;
wire na1068_2_i;
wire na1069_1;
wire na1069_1_i;
wire na1070_1;
wire na1070_1_i;
wire na1071_1;
wire na1071_1_i;
wire na1072_2;
wire na1072_2_i;
wire na1073_1;
wire na1073_1_i;
wire na1074_2;
wire na1074_2_i;
wire na1075_1;
wire na1075_1_i;
wire na1076_2;
wire na1076_2_i;
wire na1077_2;
wire na1077_2_i;
wire na1078_2;
wire na1078_2_i;
wire na1079_1;
wire na1079_1_i;
wire na1080_2;
wire na1080_2_i;
wire na1081_1;
wire na1081_1_i;
wire na1082_2;
wire na1082_2_i;
wire na1083_1;
wire na1083_1_i;
wire na1084_1;
wire na1084_1_i;
wire na1085_1;
wire na1085_1_i;
wire na1086_2;
wire na1086_2_i;
wire na1087_1;
wire na1087_1_i;
wire na1088_2;
wire na1088_2_i;
wire na1089_1;
wire na1089_1_i;
wire na1090_2;
wire na1090_2_i;
wire na1091_2;
wire na1091_2_i;
wire na1092_2;
wire na1092_2_i;
wire na1093_1;
wire na1093_1_i;
wire na1094_2;
wire na1094_2_i;
wire na1095_1;
wire na1095_1_i;
wire na1096_2;
wire na1096_2_i;
wire na1097_1;
wire na1097_1_i;
wire na1098_1;
wire na1098_1_i;
wire na1099_1;
wire na1099_1_i;
wire na1100_2;
wire na1100_2_i;
wire na1101_1;
wire na1101_1_i;
wire na1102_2;
wire na1102_2_i;
wire na1103_1;
wire na1103_1_i;
wire na1104_2;
wire na1104_2_i;
wire na1105_2;
wire na1105_2_i;
wire na1106_2;
wire na1106_2_i;
wire na1107_1;
wire na1107_1_i;
wire na1108_2;
wire na1108_2_i;
wire na1109_1;
wire na1109_1_i;
wire na1110_2;
wire na1110_2_i;
wire na1111_1;
wire na1111_1_i;
wire na1112_1;
wire na1112_1_i;
wire na1113_1;
wire na1113_1_i;
wire na1114_2;
wire na1114_2_i;
wire na1115_1;
wire na1115_1_i;
wire na1116_2;
wire na1116_2_i;
wire na1117_1;
wire na1117_1_i;
wire na1118_2;
wire na1118_2_i;
wire na1119_2;
wire na1119_2_i;
wire na1120_2;
wire na1120_2_i;
wire na1121_1;
wire na1121_1_i;
wire na1122_2;
wire na1122_2_i;
wire na1123_1;
wire na1123_1_i;
wire na1124_2;
wire na1124_2_i;
wire na1125_1;
wire na1125_1_i;
wire na1126_1;
wire na1126_1_i;
wire na1127_1;
wire na1127_1_i;
wire na1128_2;
wire na1128_2_i;
wire na1129_1;
wire na1129_1_i;
wire na1130_2;
wire na1130_2_i;
wire na1131_1;
wire na1131_1_i;
wire na1132_2;
wire na1132_2_i;
wire na1133_2;
wire na1133_2_i;
wire na1134_2;
wire na1134_2_i;
wire na1135_1;
wire na1135_1_i;
wire na1136_2;
wire na1136_2_i;
wire na1137_1;
wire na1137_1_i;
wire na1138_2;
wire na1138_2_i;
wire na1139_1;
wire na1139_1_i;
wire na1140_1;
wire na1140_1_i;
wire na1141_1;
wire na1141_1_i;
wire na1142_2;
wire na1142_2_i;
wire na1143_1;
wire na1143_1_i;
wire na1144_2;
wire na1144_2_i;
wire na1145_1;
wire na1145_1_i;
wire na1146_2;
wire na1146_2_i;
wire na1147_2;
wire na1147_2_i;
wire na1148_2;
wire na1148_2_i;
wire na1149_1;
wire na1149_1_i;
wire na1150_2;
wire na1150_2_i;
wire na1151_1;
wire na1151_1_i;
wire na1152_2;
wire na1152_2_i;
wire na1153_1;
wire na1153_1_i;
wire na1154_1;
wire na1154_1_i;
wire na1155_1;
wire na1155_1_i;
wire na1156_2;
wire na1156_2_i;
wire na1157_1;
wire na1157_1_i;
wire na1158_2;
wire na1158_2_i;
wire na1159_1;
wire na1159_1_i;
wire na1160_2;
wire na1160_2_i;
wire na1161_2;
wire na1161_2_i;
wire na1162_2;
wire na1162_2_i;
wire na1163_1;
wire na1163_1_i;
wire na1164_2;
wire na1164_2_i;
wire na1165_1;
wire na1165_1_i;
wire na1166_2;
wire na1166_2_i;
wire na1167_1;
wire na1167_1_i;
wire na1168_1;
wire na1168_1_i;
wire na1169_1;
wire na1169_1_i;
wire na1170_2;
wire na1170_2_i;
wire na1171_1;
wire na1171_1_i;
wire na1172_2;
wire na1172_2_i;
wire na1173_1;
wire na1173_1_i;
wire na1174_2;
wire na1174_2_i;
wire na1175_2;
wire na1175_2_i;
wire na1176_2;
wire na1176_2_i;
wire na1177_1;
wire na1177_1_i;
wire na1178_2;
wire na1178_2_i;
wire na1179_1;
wire na1179_1_i;
wire na1180_2;
wire na1180_2_i;
wire na1181_1;
wire na1181_1_i;
wire na1182_1;
wire na1182_1_i;
wire na1183_1;
wire na1183_1_i;
wire na1184_2;
wire na1184_2_i;
wire na1185_1;
wire na1185_1_i;
wire na1186_2;
wire na1186_2_i;
wire na1187_1;
wire na1187_1_i;
wire na1188_2;
wire na1188_2_i;
wire na1189_2;
wire na1189_2_i;
wire na1190_2;
wire na1190_2_i;
wire na1191_1;
wire na1191_1_i;
wire na1192_2;
wire na1192_2_i;
wire na1193_1;
wire na1193_1_i;
wire na1194_2;
wire na1194_2_i;
wire na1195_1;
wire na1195_1_i;
wire na1196_1;
wire na1196_1_i;
wire na1197_1;
wire na1197_1_i;
wire na1198_2;
wire na1198_2_i;
wire na1199_1;
wire na1199_1_i;
wire na1200_2;
wire na1200_2_i;
wire na1201_1;
wire na1201_1_i;
wire na1202_2;
wire na1202_2_i;
wire na1203_2;
wire na1203_2_i;
wire na1204_2;
wire na1204_2_i;
wire na1205_1;
wire na1205_1_i;
wire na1206_2;
wire na1206_2_i;
wire na1207_1;
wire na1207_1_i;
wire na1208_2;
wire na1208_2_i;
wire na1209_1;
wire na1209_1_i;
wire na1210_1;
wire na1210_1_i;
wire na1211_1;
wire na1211_1_i;
wire na1212_2;
wire na1212_2_i;
wire na1213_1;
wire na1213_1_i;
wire na1214_2;
wire na1214_2_i;
wire na1215_1;
wire na1215_1_i;
wire na1216_2;
wire na1216_2_i;
wire na1217_2;
wire na1217_2_i;
wire na1218_2;
wire na1218_2_i;
wire na1219_1;
wire na1219_1_i;
wire na1220_2;
wire na1220_2_i;
wire na1221_1;
wire na1221_1_i;
wire na1222_2;
wire na1222_2_i;
wire na1223_1;
wire na1223_1_i;
wire na1224_1;
wire na1224_1_i;
wire na1225_1;
wire na1225_1_i;
wire na1226_2;
wire na1226_2_i;
wire na1227_1;
wire na1227_1_i;
wire na1228_2;
wire na1228_2_i;
wire na1229_1;
wire na1229_1_i;
wire na1230_2;
wire na1230_2_i;
wire na1231_2;
wire na1231_2_i;
wire na1232_2;
wire na1232_2_i;
wire na1233_1;
wire na1233_1_i;
wire na1234_2;
wire na1234_2_i;
wire na1235_1;
wire na1235_1_i;
wire na1236_2;
wire na1236_2_i;
wire na1237_1;
wire na1237_1_i;
wire na1238_1;
wire na1238_1_i;
wire na1239_1;
wire na1239_1_i;
wire na1240_2;
wire na1240_2_i;
wire na1241_1;
wire na1241_1_i;
wire na1242_2;
wire na1242_2_i;
wire na1243_1;
wire na1243_1_i;
wire na1244_2;
wire na1244_2_i;
wire na1245_2;
wire na1245_2_i;
wire na1246_2;
wire na1246_2_i;
wire na1247_1;
wire na1247_1_i;
wire na1248_2;
wire na1248_2_i;
wire na1249_1;
wire na1249_1_i;
wire na1250_2;
wire na1250_2_i;
wire na1251_1;
wire na1251_1_i;
wire na1252_1;
wire na1252_1_i;
wire na1253_1;
wire na1253_1_i;
wire na1254_2;
wire na1254_2_i;
wire na1255_1;
wire na1255_1_i;
wire na1256_2;
wire na1256_2_i;
wire na1257_1;
wire na1257_1_i;
wire na1258_2;
wire na1258_2_i;
wire na1259_2;
wire na1259_2_i;
wire na1260_2;
wire na1260_2_i;
wire na1261_1;
wire na1261_1_i;
wire na1262_2;
wire na1262_2_i;
wire na1263_1;
wire na1263_1_i;
wire na1264_2;
wire na1264_2_i;
wire na1265_1;
wire na1265_1_i;
wire na1266_1;
wire na1266_1_i;
wire na1267_1;
wire na1267_1_i;
wire na1268_2;
wire na1268_2_i;
wire na1269_1;
wire na1269_1_i;
wire na1270_2;
wire na1270_2_i;
wire na1271_1;
wire na1271_1_i;
wire na1272_2;
wire na1272_2_i;
wire na1273_2;
wire na1273_2_i;
wire na1274_2;
wire na1274_2_i;
wire na1275_1;
wire na1275_1_i;
wire na1276_2;
wire na1276_2_i;
wire na1277_1;
wire na1277_1_i;
wire na1278_2;
wire na1278_2_i;
wire na1279_1;
wire na1279_1_i;
wire na1280_1;
wire na1280_1_i;
wire na1281_1;
wire na1281_1_i;
wire na1282_2;
wire na1282_2_i;
wire na1283_1;
wire na1283_1_i;
wire na1284_2;
wire na1284_2_i;
wire na1285_1;
wire na1285_1_i;
wire na1286_2;
wire na1286_2_i;
wire na1287_2;
wire na1287_2_i;
wire na1288_2;
wire na1288_2_i;
wire na1289_1;
wire na1289_1_i;
wire na1290_2;
wire na1290_2_i;
wire na1291_1;
wire na1291_1_i;
wire na1292_2;
wire na1292_2_i;
wire na1293_1;
wire na1293_1_i;
wire na1294_1;
wire na1294_1_i;
wire na1295_1;
wire na1295_1_i;
wire na1296_2;
wire na1296_2_i;
wire na1297_1;
wire na1297_1_i;
wire na1298_2;
wire na1298_2_i;
wire na1299_1;
wire na1299_1_i;
wire na1300_2;
wire na1300_2_i;
wire na1301_2;
wire na1301_2_i;
wire na1302_2;
wire na1302_2_i;
wire na1303_1;
wire na1303_1_i;
wire na1304_2;
wire na1304_2_i;
wire na1305_1;
wire na1305_1_i;
wire na1306_2;
wire na1306_2_i;
wire na1307_1;
wire na1307_1_i;
wire na1308_1;
wire na1308_1_i;
wire na1309_1;
wire na1309_1_i;
wire na1310_2;
wire na1310_2_i;
wire na1311_1;
wire na1311_1_i;
wire na1312_2;
wire na1312_2_i;
wire na1313_1;
wire na1313_1_i;
wire na1314_2;
wire na1314_2_i;
wire na1315_2;
wire na1315_2_i;
wire na1316_2;
wire na1316_2_i;
wire na1317_1;
wire na1317_1_i;
wire na1318_2;
wire na1318_2_i;
wire na1319_1;
wire na1319_1_i;
wire na1320_2;
wire na1320_2_i;
wire na1321_1;
wire na1321_1_i;
wire na1322_1;
wire na1322_1_i;
wire na1323_1;
wire na1323_1_i;
wire na1324_2;
wire na1324_2_i;
wire na1325_1;
wire na1325_1_i;
wire na1326_2;
wire na1326_2_i;
wire na1327_1;
wire na1327_1_i;
wire na1328_2;
wire na1328_2_i;
wire na1329_2;
wire na1329_2_i;
wire na1330_2;
wire na1330_2_i;
wire na1331_1;
wire na1331_1_i;
wire na1332_2;
wire na1332_2_i;
wire na1333_1;
wire na1333_1_i;
wire na1334_2;
wire na1334_2_i;
wire na1335_1;
wire na1335_1_i;
wire na1336_1;
wire na1336_1_i;
wire na1337_1;
wire na1337_1_i;
wire na1338_2;
wire na1338_2_i;
wire na1339_1;
wire na1339_1_i;
wire na1340_2;
wire na1340_2_i;
wire na1341_1;
wire na1341_1_i;
wire na1342_2;
wire na1342_2_i;
wire na1343_2;
wire na1343_2_i;
wire na1344_2;
wire na1344_2_i;
wire na1345_1;
wire na1345_1_i;
wire na1346_2;
wire na1346_2_i;
wire na1347_1;
wire na1347_1_i;
wire na1348_2;
wire na1348_2_i;
wire na1349_1;
wire na1349_1_i;
wire na1350_1;
wire na1350_1_i;
wire na1351_1;
wire na1351_1_i;
wire na1352_2;
wire na1352_2_i;
wire na1353_1;
wire na1353_1_i;
wire na1354_2;
wire na1354_2_i;
wire na1355_1;
wire na1355_1_i;
wire na1356_2;
wire na1356_2_i;
wire na1357_2;
wire na1357_2_i;
wire na1358_2;
wire na1358_2_i;
wire na1359_1;
wire na1359_1_i;
wire na1360_2;
wire na1360_2_i;
wire na1361_1;
wire na1361_1_i;
wire na1362_2;
wire na1362_2_i;
wire na1363_1;
wire na1363_1_i;
wire na1364_1;
wire na1364_1_i;
wire na1365_1;
wire na1365_1_i;
wire na1366_2;
wire na1366_2_i;
wire na1367_1;
wire na1367_1_i;
wire na1368_2;
wire na1368_2_i;
wire na1369_1;
wire na1369_1_i;
wire na1370_2;
wire na1370_2_i;
wire na1371_2;
wire na1371_2_i;
wire na1372_2;
wire na1372_2_i;
wire na1373_1;
wire na1373_1_i;
wire na1374_2;
wire na1374_2_i;
wire na1375_1;
wire na1375_1_i;
wire na1376_2;
wire na1376_2_i;
wire na1377_1;
wire na1377_1_i;
wire na1378_1;
wire na1378_1_i;
wire na1379_1;
wire na1379_1_i;
wire na1380_2;
wire na1380_2_i;
wire na1381_1;
wire na1381_1_i;
wire na1382_2;
wire na1382_2_i;
wire na1383_1;
wire na1383_1_i;
wire na1384_2;
wire na1384_2_i;
wire na1385_2;
wire na1385_2_i;
wire na1386_2;
wire na1386_2_i;
wire na1387_1;
wire na1387_1_i;
wire na1388_2;
wire na1388_2_i;
wire na1389_1;
wire na1389_1_i;
wire na1390_2;
wire na1390_2_i;
wire na1391_1;
wire na1391_1_i;
wire na1392_1;
wire na1392_1_i;
wire na1393_1;
wire na1393_1_i;
wire na1394_2;
wire na1394_2_i;
wire na1395_1;
wire na1395_1_i;
wire na1396_2;
wire na1396_2_i;
wire na1397_1;
wire na1397_1_i;
wire na1398_2;
wire na1398_2_i;
wire na1399_2;
wire na1399_2_i;
wire na1400_2;
wire na1400_2_i;
wire na1401_1;
wire na1401_1_i;
wire na1402_2;
wire na1402_2_i;
wire na1403_1;
wire na1403_1_i;
wire na1404_2;
wire na1404_2_i;
wire na1405_1;
wire na1405_1_i;
wire na1406_1;
wire na1406_1_i;
wire na1407_1;
wire na1407_1_i;
wire na1408_2;
wire na1408_2_i;
wire na1409_1;
wire na1409_1_i;
wire na1410_2;
wire na1410_2_i;
wire na1411_1;
wire na1411_1_i;
wire na1412_2;
wire na1412_2_i;
wire na1413_2;
wire na1413_2_i;
wire na1414_2;
wire na1414_2_i;
wire na1415_1;
wire na1415_1_i;
wire na1416_2;
wire na1416_2_i;
wire na1417_1;
wire na1417_1_i;
wire na1418_2;
wire na1418_2_i;
wire na1419_1;
wire na1419_1_i;
wire na1420_1;
wire na1420_1_i;
wire na1421_1;
wire na1421_1_i;
wire na1422_2;
wire na1422_2_i;
wire na1423_1;
wire na1423_1_i;
wire na1424_2;
wire na1424_2_i;
wire na1425_1;
wire na1425_1_i;
wire na1426_2;
wire na1426_2_i;
wire na1427_2;
wire na1427_2_i;
wire na1428_2;
wire na1428_2_i;
wire na1429_1;
wire na1429_1_i;
wire na1430_2;
wire na1430_2_i;
wire na1431_1;
wire na1431_1_i;
wire na1432_2;
wire na1432_2_i;
wire na1433_1;
wire na1433_1_i;
wire na1434_1;
wire na1434_1_i;
wire na1435_1;
wire na1435_1_i;
wire na1436_2;
wire na1436_2_i;
wire na1437_1;
wire na1437_1_i;
wire na1438_2;
wire na1438_2_i;
wire na1439_1;
wire na1439_1_i;
wire na1440_2;
wire na1440_2_i;
wire na1441_2;
wire na1441_2_i;
wire na1442_2;
wire na1442_2_i;
wire na1443_1;
wire na1443_1_i;
wire na1444_2;
wire na1444_2_i;
wire na1445_1;
wire na1445_1_i;
wire na1446_2;
wire na1446_2_i;
wire na1447_1;
wire na1447_1_i;
wire na1448_1;
wire na1448_1_i;
wire na1449_1;
wire na1449_1_i;
wire na1450_2;
wire na1450_2_i;
wire na1451_1;
wire na1451_1_i;
wire na1452_2;
wire na1452_2_i;
wire na1453_1;
wire na1453_1_i;
wire na1454_2;
wire na1454_2_i;
wire na1455_2;
wire na1455_2_i;
wire na1456_2;
wire na1456_2_i;
wire na1457_1;
wire na1457_1_i;
wire na1458_2;
wire na1458_2_i;
wire na1459_1;
wire na1459_1_i;
wire na1460_2;
wire na1460_2_i;
wire na1461_1;
wire na1461_1_i;
wire na1462_1;
wire na1462_1_i;
wire na1463_1;
wire na1463_1_i;
wire na1464_2;
wire na1464_2_i;
wire na1465_1;
wire na1465_1_i;
wire na1466_2;
wire na1466_2_i;
wire na1467_1;
wire na1467_1_i;
wire na1468_2;
wire na1468_2_i;
wire na1469_2;
wire na1469_2_i;
wire na1470_2;
wire na1470_2_i;
wire na1471_1;
wire na1471_1_i;
wire na1472_2;
wire na1472_2_i;
wire na1473_1;
wire na1473_1_i;
wire na1474_2;
wire na1474_2_i;
wire na1475_1;
wire na1475_1_i;
wire na1476_1;
wire na1476_1_i;
wire na1477_1;
wire na1477_1_i;
wire na1478_2;
wire na1478_2_i;
wire na1479_1;
wire na1479_1_i;
wire na1480_2;
wire na1480_2_i;
wire na1481_1;
wire na1481_1_i;
wire na1482_2;
wire na1482_2_i;
wire na1483_2;
wire na1483_2_i;
wire na1484_2;
wire na1484_2_i;
wire na1485_1;
wire na1485_1_i;
wire na1486_2;
wire na1486_2_i;
wire na1487_1;
wire na1487_1_i;
wire na1488_2;
wire na1488_2_i;
wire na1489_1;
wire na1489_1_i;
wire na1490_1;
wire na1490_1_i;
wire na1491_1;
wire na1491_1_i;
wire na1492_2;
wire na1492_2_i;
wire na1493_1;
wire na1493_1_i;
wire na1494_2;
wire na1494_2_i;
wire na1495_1;
wire na1495_1_i;
wire na1496_2;
wire na1496_2_i;
wire na1497_2;
wire na1497_2_i;
wire na1498_2;
wire na1498_2_i;
wire na1499_1;
wire na1499_1_i;
wire na1500_2;
wire na1500_2_i;
wire na1501_1;
wire na1501_1_i;
wire na1502_2;
wire na1502_2_i;
wire na1503_1;
wire na1503_1_i;
wire na1504_1;
wire na1504_1_i;
wire na1505_1;
wire na1505_1_i;
wire na1506_2;
wire na1506_2_i;
wire na1507_1;
wire na1507_1_i;
wire na1508_2;
wire na1508_2_i;
wire na1509_1;
wire na1509_1_i;
wire na1510_2;
wire na1510_2_i;
wire na1511_2;
wire na1511_2_i;
wire na1512_2;
wire na1512_2_i;
wire na1513_1;
wire na1513_1_i;
wire na1514_2;
wire na1514_2_i;
wire na1515_1;
wire na1515_1_i;
wire na1516_2;
wire na1516_2_i;
wire na1517_1;
wire na1517_1_i;
wire na1518_1;
wire na1518_1_i;
wire na1519_1;
wire na1519_1_i;
wire na1520_2;
wire na1520_2_i;
wire na1521_1;
wire na1521_1_i;
wire na1522_2;
wire na1522_2_i;
wire na1523_1;
wire na1523_1_i;
wire na1524_2;
wire na1524_2_i;
wire na1525_2;
wire na1525_2_i;
wire na1526_2;
wire na1526_2_i;
wire na1527_1;
wire na1527_1_i;
wire na1528_2;
wire na1528_2_i;
wire na1529_1;
wire na1529_1_i;
wire na1530_2;
wire na1530_2_i;
wire na1531_1;
wire na1531_1_i;
wire na1532_1;
wire na1532_1_i;
wire na1533_1;
wire na1533_1_i;
wire na1534_2;
wire na1534_2_i;
wire na1535_1;
wire na1535_1_i;
wire na1536_2;
wire na1536_2_i;
wire na1537_1;
wire na1537_1_i;
wire na1538_2;
wire na1538_2_i;
wire na1539_2;
wire na1539_2_i;
wire na1540_2;
wire na1540_2_i;
wire na1541_1;
wire na1541_1_i;
wire na1542_2;
wire na1542_2_i;
wire na1543_1;
wire na1543_1_i;
wire na1544_2;
wire na1544_2_i;
wire na1545_1;
wire na1545_1_i;
wire na1546_1;
wire na1546_1_i;
wire na1547_1;
wire na1547_1_i;
wire na1548_2;
wire na1548_2_i;
wire na1549_1;
wire na1549_1_i;
wire na1550_2;
wire na1550_2_i;
wire na1551_1;
wire na1551_1_i;
wire na1552_2;
wire na1552_2_i;
wire na1553_2;
wire na1553_2_i;
wire na1554_2;
wire na1554_2_i;
wire na1555_1;
wire na1555_1_i;
wire na1556_2;
wire na1556_2_i;
wire na1557_1;
wire na1557_1_i;
wire na1558_2;
wire na1558_2_i;
wire na1559_1;
wire na1559_1_i;
wire na1560_1;
wire na1560_1_i;
wire na1561_1;
wire na1561_1_i;
wire na1562_2;
wire na1562_2_i;
wire na1563_1;
wire na1563_1_i;
wire na1564_2;
wire na1564_2_i;
wire na1565_1;
wire na1565_1_i;
wire na1566_2;
wire na1566_2_i;
wire na1567_2;
wire na1567_2_i;
wire na1568_2;
wire na1568_2_i;
wire na1569_1;
wire na1569_1_i;
wire na1570_2;
wire na1570_2_i;
wire na1571_1;
wire na1571_1_i;
wire na1572_2;
wire na1572_2_i;
wire na1573_1;
wire na1573_1_i;
wire na1574_1;
wire na1574_1_i;
wire na1575_1;
wire na1575_1_i;
wire na1576_2;
wire na1576_2_i;
wire na1577_1;
wire na1577_1_i;
wire na1578_2;
wire na1578_2_i;
wire na1579_1;
wire na1579_1_i;
wire na1580_2;
wire na1580_2_i;
wire na1581_2;
wire na1581_2_i;
wire na1582_2;
wire na1582_2_i;
wire na1583_1;
wire na1583_1_i;
wire na1584_2;
wire na1584_2_i;
wire na1585_1;
wire na1585_1_i;
wire na1586_2;
wire na1586_2_i;
wire na1587_1;
wire na1587_1_i;
wire na1588_1;
wire na1588_1_i;
wire na1589_1;
wire na1589_1_i;
wire na1590_2;
wire na1590_2_i;
wire na1591_1;
wire na1591_1_i;
wire na1592_2;
wire na1592_2_i;
wire na1593_1;
wire na1593_1_i;
wire na1594_2;
wire na1594_2_i;
wire na1595_2;
wire na1595_2_i;
wire na1596_2;
wire na1596_2_i;
wire na1597_1;
wire na1597_1_i;
wire na1598_2;
wire na1598_2_i;
wire na1599_1;
wire na1599_1_i;
wire na1600_2;
wire na1600_2_i;
wire na1601_1;
wire na1601_1_i;
wire na1602_1;
wire na1602_1_i;
wire na1603_1;
wire na1603_1_i;
wire na1604_2;
wire na1604_2_i;
wire na1605_1;
wire na1605_1_i;
wire na1606_2;
wire na1606_2_i;
wire na1607_1;
wire na1607_1_i;
wire na1608_2;
wire na1608_2_i;
wire na1609_2;
wire na1609_2_i;
wire na1610_2;
wire na1610_2_i;
wire na1611_1;
wire na1611_1_i;
wire na1612_2;
wire na1612_2_i;
wire na1613_1;
wire na1613_1_i;
wire na1614_2;
wire na1614_2_i;
wire na1615_1;
wire na1615_1_i;
wire na1616_1;
wire na1616_1_i;
wire na1617_1;
wire na1617_1_i;
wire na1618_2;
wire na1618_2_i;
wire na1619_1;
wire na1619_1_i;
wire na1620_2;
wire na1620_2_i;
wire na1621_1;
wire na1621_1_i;
wire na1622_2;
wire na1622_2_i;
wire na1623_2;
wire na1623_2_i;
wire na1624_2;
wire na1624_2_i;
wire na1625_1;
wire na1625_1_i;
wire na1626_2;
wire na1626_2_i;
wire na1627_1;
wire na1627_1_i;
wire na1628_2;
wire na1628_2_i;
wire na1629_1;
wire na1629_1_i;
wire na1630_1;
wire na1630_1_i;
wire na1631_1;
wire na1631_1_i;
wire na1632_2;
wire na1632_2_i;
wire na1633_1;
wire na1633_1_i;
wire na1634_2;
wire na1634_2_i;
wire na1635_1;
wire na1635_1_i;
wire na1636_2;
wire na1636_2_i;
wire na1637_2;
wire na1637_2_i;
wire na1638_2;
wire na1638_2_i;
wire na1639_1;
wire na1639_1_i;
wire na1640_2;
wire na1640_2_i;
wire na1641_1;
wire na1641_1_i;
wire na1642_2;
wire na1642_2_i;
wire na1643_1;
wire na1643_1_i;
wire na1644_1;
wire na1644_1_i;
wire na1645_1;
wire na1645_1_i;
wire na1646_2;
wire na1646_2_i;
wire na1647_1;
wire na1647_1_i;
wire na1648_2;
wire na1648_2_i;
wire na1649_1;
wire na1649_1_i;
wire na1650_2;
wire na1650_2_i;
wire na1651_2;
wire na1651_2_i;
wire na1652_2;
wire na1652_2_i;
wire na1653_1;
wire na1653_1_i;
wire na1654_2;
wire na1654_2_i;
wire na1655_1;
wire na1655_1_i;
wire na1656_2;
wire na1656_2_i;
wire na1657_1;
wire na1657_1_i;
wire na1658_1;
wire na1658_1_i;
wire na1659_1;
wire na1659_1_i;
wire na1660_2;
wire na1660_2_i;
wire na1661_1;
wire na1661_1_i;
wire na1662_2;
wire na1662_2_i;
wire na1663_1;
wire na1663_1_i;
wire na1664_2;
wire na1664_2_i;
wire na1665_2;
wire na1665_2_i;
wire na1666_2;
wire na1666_2_i;
wire na1667_1;
wire na1667_1_i;
wire na1668_2;
wire na1668_2_i;
wire na1669_1;
wire na1669_1_i;
wire na1670_2;
wire na1670_2_i;
wire na1671_1;
wire na1671_1_i;
wire na1672_1;
wire na1672_1_i;
wire na1673_1;
wire na1673_1_i;
wire na1674_2;
wire na1674_2_i;
wire na1675_1;
wire na1675_1_i;
wire na1676_2;
wire na1676_2_i;
wire na1677_1;
wire na1677_1_i;
wire na1678_2;
wire na1678_2_i;
wire na1679_2;
wire na1679_2_i;
wire na1680_2;
wire na1680_2_i;
wire na1681_1;
wire na1681_1_i;
wire na1682_2;
wire na1682_2_i;
wire na1683_1;
wire na1683_1_i;
wire na1684_2;
wire na1684_2_i;
wire na1685_1;
wire na1685_1_i;
wire na1686_1;
wire na1686_1_i;
wire na1687_1;
wire na1687_1_i;
wire na1688_2;
wire na1688_2_i;
wire na1689_1;
wire na1689_1_i;
wire na1690_2;
wire na1690_2_i;
wire na1691_1;
wire na1691_1_i;
wire na1692_2;
wire na1692_2_i;
wire na1693_2;
wire na1693_2_i;
wire na1694_2;
wire na1694_2_i;
wire na1695_1;
wire na1695_1_i;
wire na1696_2;
wire na1696_2_i;
wire na1697_1;
wire na1697_1_i;
wire na1698_2;
wire na1698_2_i;
wire na1699_1;
wire na1699_1_i;
wire na1700_1;
wire na1700_1_i;
wire na1701_1;
wire na1701_1_i;
wire na1702_2;
wire na1702_2_i;
wire na1703_1;
wire na1703_1_i;
wire na1704_2;
wire na1704_2_i;
wire na1705_1;
wire na1705_1_i;
wire na1706_2;
wire na1706_2_i;
wire na1707_2;
wire na1707_2_i;
wire na1708_2;
wire na1708_2_i;
wire na1709_1;
wire na1709_1_i;
wire na1710_2;
wire na1710_2_i;
wire na1711_1;
wire na1711_1_i;
wire na1712_2;
wire na1712_2_i;
wire na1713_1;
wire na1713_1_i;
wire na1714_1;
wire na1714_1_i;
wire na1715_1;
wire na1715_1_i;
wire na1716_2;
wire na1716_2_i;
wire na1717_1;
wire na1717_1_i;
wire na1718_2;
wire na1718_2_i;
wire na1719_1;
wire na1719_1_i;
wire na1720_2;
wire na1720_2_i;
wire na1721_2;
wire na1721_2_i;
wire na1722_2;
wire na1722_2_i;
wire na1723_1;
wire na1723_1_i;
wire na1724_2;
wire na1724_2_i;
wire na1725_1;
wire na1725_1_i;
wire na1726_2;
wire na1726_2_i;
wire na1727_1;
wire na1727_1_i;
wire na1728_1;
wire na1728_1_i;
wire na1729_1;
wire na1729_1_i;
wire na1730_2;
wire na1730_2_i;
wire na1731_1;
wire na1731_1_i;
wire na1732_2;
wire na1732_2_i;
wire na1733_1;
wire na1733_1_i;
wire na1734_2;
wire na1734_2_i;
wire na1735_2;
wire na1735_2_i;
wire na1736_2;
wire na1736_2_i;
wire na1737_1;
wire na1737_1_i;
wire na1738_2;
wire na1738_2_i;
wire na1739_1;
wire na1739_1_i;
wire na1740_2;
wire na1740_2_i;
wire na1741_1;
wire na1741_1_i;
wire na1742_1;
wire na1742_1_i;
wire na1743_1;
wire na1743_1_i;
wire na1744_2;
wire na1744_2_i;
wire na1745_1;
wire na1745_1_i;
wire na1746_2;
wire na1746_2_i;
wire na1747_1;
wire na1747_1_i;
wire na1748_2;
wire na1748_2_i;
wire na1749_2;
wire na1749_2_i;
wire na1750_2;
wire na1750_2_i;
wire na1751_1;
wire na1751_1_i;
wire na1752_2;
wire na1752_2_i;
wire na1753_1;
wire na1753_1_i;
wire na1754_2;
wire na1754_2_i;
wire na1755_1;
wire na1755_1_i;
wire na1756_1;
wire na1756_1_i;
wire na1757_1;
wire na1757_1_i;
wire na1758_2;
wire na1758_2_i;
wire na1759_1;
wire na1759_1_i;
wire na1760_2;
wire na1760_2_i;
wire na1761_1;
wire na1761_1_i;
wire na1762_2;
wire na1762_2_i;
wire na1763_2;
wire na1763_2_i;
wire na1764_2;
wire na1764_2_i;
wire na1765_1;
wire na1765_1_i;
wire na1766_2;
wire na1766_2_i;
wire na1767_1;
wire na1767_1_i;
wire na1768_2;
wire na1768_2_i;
wire na1769_1;
wire na1769_1_i;
wire na1770_1;
wire na1770_1_i;
wire na1771_1;
wire na1771_1_i;
wire na1772_2;
wire na1772_2_i;
wire na1773_1;
wire na1773_1_i;
wire na1774_2;
wire na1774_2_i;
wire na1775_1;
wire na1775_1_i;
wire na1776_2;
wire na1776_2_i;
wire na1777_2;
wire na1777_2_i;
wire na1778_2;
wire na1778_2_i;
wire na1779_1;
wire na1779_1_i;
wire na1780_2;
wire na1780_2_i;
wire na1781_1;
wire na1781_1_i;
wire na1782_2;
wire na1782_2_i;
wire na1783_1;
wire na1783_1_i;
wire na1784_1;
wire na1784_1_i;
wire na1785_1;
wire na1785_1_i;
wire na1786_2;
wire na1786_2_i;
wire na1787_1;
wire na1787_1_i;
wire na1788_2;
wire na1788_2_i;
wire na1789_1;
wire na1789_1_i;
wire na1790_2;
wire na1790_2_i;
wire na1791_2;
wire na1791_2_i;
wire na1792_2;
wire na1792_2_i;
wire na1793_1;
wire na1793_1_i;
wire na1794_2;
wire na1794_2_i;
wire na1795_1;
wire na1795_1_i;
wire na1796_2;
wire na1796_2_i;
wire na1797_1;
wire na1797_1_i;
wire na1798_1;
wire na1798_1_i;
wire na1799_1;
wire na1799_1_i;
wire na1800_2;
wire na1800_2_i;
wire na1801_1;
wire na1801_1_i;
wire na1802_2;
wire na1802_2_i;
wire na1803_1;
wire na1803_1_i;
wire na1804_2;
wire na1804_2_i;
wire na1805_2;
wire na1805_2_i;
wire na1806_2;
wire na1806_2_i;
wire na1807_1;
wire na1807_1_i;
wire na1808_2;
wire na1808_2_i;
wire na1809_1;
wire na1809_1_i;
wire na1810_2;
wire na1810_2_i;
wire na1811_1;
wire na1811_1_i;
wire na1812_1;
wire na1812_1_i;
wire na1813_1;
wire na1813_1_i;
wire na1814_2;
wire na1814_2_i;
wire na1815_1;
wire na1815_1_i;
wire na1816_2;
wire na1816_2_i;
wire na1817_1;
wire na1817_1_i;
wire na1818_2;
wire na1818_2_i;
wire na1819_2;
wire na1819_2_i;
wire na1820_2;
wire na1820_2_i;
wire na1821_1;
wire na1821_1_i;
wire na1822_2;
wire na1822_2_i;
wire na1823_1;
wire na1823_1_i;
wire na1824_2;
wire na1824_2_i;
wire na1825_1;
wire na1825_1_i;
wire na1826_1;
wire na1826_1_i;
wire na1827_1;
wire na1827_1_i;
wire na1828_2;
wire na1828_2_i;
wire na1829_1;
wire na1829_1_i;
wire na1830_2;
wire na1830_2_i;
wire na1831_1;
wire na1831_1_i;
wire na1832_2;
wire na1832_2_i;
wire na1833_2;
wire na1833_2_i;
wire na1834_2;
wire na1834_2_i;
wire na1835_1;
wire na1835_1_i;
wire na1836_2;
wire na1836_2_i;
wire na1837_1;
wire na1837_1_i;
wire na1838_2;
wire na1838_2_i;
wire na1839_1;
wire na1839_1_i;
wire na1840_1;
wire na1840_1_i;
wire na1841_1;
wire na1841_1_i;
wire na1842_2;
wire na1842_2_i;
wire na1843_1;
wire na1843_1_i;
wire na1844_2;
wire na1844_2_i;
wire na1845_1;
wire na1845_1_i;
wire na1846_2;
wire na1846_2_i;
wire na1847_2;
wire na1847_2_i;
wire na1848_2;
wire na1848_2_i;
wire na1849_1;
wire na1849_1_i;
wire na1850_2;
wire na1850_2_i;
wire na1851_1;
wire na1851_1_i;
wire na1852_2;
wire na1852_2_i;
wire na1853_1;
wire na1853_1_i;
wire na1854_1;
wire na1854_1_i;
wire na1855_1;
wire na1855_1_i;
wire na1856_2;
wire na1856_2_i;
wire na1857_1;
wire na1857_1_i;
wire na1858_2;
wire na1858_2_i;
wire na1859_1;
wire na1859_1_i;
wire na1860_2;
wire na1860_2_i;
wire na1861_2;
wire na1861_2_i;
wire na1862_2;
wire na1862_2_i;
wire na1863_1;
wire na1863_1_i;
wire na1864_2;
wire na1864_2_i;
wire na1865_1;
wire na1865_1_i;
wire na1866_2;
wire na1866_2_i;
wire na1867_1;
wire na1867_1_i;
wire na1868_1;
wire na1868_1_i;
wire na1869_1;
wire na1869_1_i;
wire na1870_2;
wire na1870_2_i;
wire na1871_1;
wire na1871_1_i;
wire na1872_2;
wire na1872_2_i;
wire na1873_1;
wire na1873_1_i;
wire na1874_2;
wire na1874_2_i;
wire na1875_2;
wire na1875_2_i;
wire na1876_2;
wire na1876_2_i;
wire na1877_1;
wire na1877_1_i;
wire na1878_2;
wire na1878_2_i;
wire na1879_1;
wire na1879_1_i;
wire na1880_2;
wire na1880_2_i;
wire na1881_1;
wire na1881_1_i;
wire na1882_1;
wire na1883_1;
wire na1884_1;
wire na1885_1;
wire na1886_1;
wire na1887_1;
wire na1888_1;
wire na1889_1;
wire na1890_1;
wire na1891_1;
wire na1892_1;
wire na1893_1;
wire na1894_1;
wire na1895_1;
wire na1896_1;
wire na1897_1;
wire na1898_1;
wire na1899_1;
wire na1900_1;
wire na1901_1;
wire na1902_1;
wire na1903_1;
wire na1904_1;
wire na1905_1;
wire na1906_1;
wire na1907_1;
wire na1908_1;
wire na1909_1;
wire na1910_1;
wire na1911_1;
wire na1912_1;
wire na1913_1;
wire na1914_1;
wire na1915_1;
wire na1916_1;
wire na1917_1;
wire na1918_1;
wire na1919_1;
wire na1920_1;
wire na1921_1;
wire na1922_1;
wire na1923_1;
wire na1924_1;
wire na1925_1;
wire na1926_1;
wire na1927_1;
wire na1928_1;
wire na1929_1;
wire na1930_1;
wire na1931_1;
wire na1932_1;
wire na1933_1;
wire na1934_1;
wire na1935_1;
wire na1936_1;
wire na1937_1;
wire na1938_1;
wire na1939_1;
wire na1940_1;
wire na1941_1;
wire na1942_1;
wire na1943_1;
wire na1944_1;
wire na1945_1;
wire na1946_1;
wire na1947_1;
wire na1948_1;
wire na1949_1;
wire na1950_1;
wire na1951_1;
wire na1952_1;
wire na1953_1;
wire na1954_1;
wire na1955_1;
wire na1956_1;
wire na1957_1;
wire na1958_1;
wire na1959_1;
wire na1960_1;
wire na1961_1;
wire na1962_1;
wire na1963_1;
wire na1964_1;
wire na1965_1;
wire na1966_1;
wire na1967_1;
wire na1968_1;
wire na1969_1;
wire na1970_1;
wire na1971_1;
wire na1972_1;
wire na1973_1;
wire na1974_1;
wire na1975_1;
wire na1976_1;
wire na1977_1;
wire na1978_1;
wire na1979_1;
wire na1980_1;
wire na1981_1;
wire na1982_1;
wire na1983_1;
wire na1984_1;
wire na1985_1;
wire na1986_1;
wire na1987_1;
wire na1988_1;
wire na1989_1;
wire na1990_1;
wire na1991_1;
wire na1992_1;
wire na1993_1;
wire na1994_1;
wire na1995_1;
wire na1996_1;
wire na1997_1;
wire na1998_1;
wire na1999_1;
wire na2000_1;
wire na2001_1;
wire na2002_1;
wire na2003_1;
wire na2004_1;
wire na2005_1;
wire na2006_1;
wire na2007_1;
wire na2008_1;
wire na2009_1;
wire na2010_1;
wire na2011_1;
wire na2012_1;
wire na2013_1;
wire na2014_1;
wire na2015_1;
wire na2016_1;
wire na2017_1;
wire na2018_1;
wire na2019_1;
wire na2020_1;
wire na2021_1;
wire na2022_1;
wire na2023_1;
wire na2024_1;
wire na2025_1;
wire na2026_1;
wire na2027_1;
wire na2028_1;
wire na2029_1;
wire na2030_1;
wire na2031_1;
wire na2032_1;
wire na2033_1;
wire na2034_1;
wire na2035_1;
wire na2036_1;
wire na2037_1;
wire na2038_1;
wire na2039_1;
wire na2040_1;
wire na2041_1;
wire na2042_1;
wire na2043_1;
wire na2044_1;
wire na2045_1;
wire na2046_1;
wire na2047_1;
wire na2048_1;
wire na2049_1;
wire na2050_1;
wire na2051_1;
wire na2052_1;
wire na2053_1;
wire na2054_1;
wire na2055_1;
wire na2056_1;
wire na2057_1;
wire na2058_1;
wire na2059_1;
wire na2060_1;
wire na2061_1;
wire na2062_1;
wire na2063_1;
wire na2064_1;
wire na2065_1;
wire na2066_1;
wire na2067_1;
wire na2068_1;
wire na2069_1;
wire na2070_1;
wire na2071_1;
wire na2072_1;
wire na2073_1;
wire na2074_1;
wire na2075_1;
wire na2076_1;
wire na2077_1;
wire na2078_1;
wire na2079_1;
wire na2080_1;
wire na2081_1;
wire na2082_1;
wire na2083_1;
wire na2084_1;
wire na2085_1;
wire na2086_1;
wire na2087_1;
wire na2088_1;
wire na2089_1;
wire na2090_1;
wire na2091_1;
wire na2092_1;
wire na2093_1;
wire na2094_1;
wire na2095_1;
wire na2096_1;
wire na2097_1;
wire na2098_1;
wire na2099_1;
wire na2100_1;
wire na2101_1;
wire na2102_1;
wire na2103_1;
wire na2104_1;
wire na2105_1;
wire na2106_1;
wire na2107_1;
wire na2108_1;
wire na2109_1;
wire na2110_1;
wire na2111_1;
wire na2112_1;
wire na2113_1;
wire na2114_1;
wire na2115_1;
wire na2116_1;
wire na2117_1;
wire na2118_1;
wire na2119_1;
wire na2120_1;
wire na2121_1;
wire na2122_1;
wire na2123_1;
wire na2124_1;
wire na2125_1;
wire na2126_1;
wire na2127_1;
wire na2128_1;
wire na2129_1;
wire na2130_1;
wire na2131_1;
wire na2132_1;
wire na2133_1;
wire na2134_1;
wire na2135_1;
wire na2136_1;
wire na2137_1;
wire na2138_1;
wire na2139_1;
wire na2140_1;
wire na2141_1;
wire na2142_1;
wire na2143_1;
wire na2144_1;
wire na2145_1;
wire na2146_1;
wire na2147_1;
wire na2148_1;
wire na2149_1;
wire na2150_1;
wire na2151_1;
wire na2152_1;
wire na2153_1;
wire na2154_1;
wire na2155_1;
wire na2156_1;
wire na2157_1;
wire na2158_1;
wire na2159_1;
wire na2160_1;
wire na2161_1;
wire na2162_1;
wire na2163_1;
wire na2164_1;
wire na2165_1;
wire na2166_1;
wire na2167_1;
wire na2168_1;
wire na2169_1;
wire na2170_1;
wire na2171_1;
wire na2172_1;
wire na2173_1;
wire na2174_1;
wire na2175_1;
wire na2176_1;
wire na2177_1;
wire na2178_1;
wire na2179_1;
wire na2180_1;
wire na2181_1;
wire na2182_1;
wire na2183_1;
wire na2184_1;
wire na2185_1;
wire na2186_1;
wire na2187_1;
wire na2188_1;
wire na2189_1;
wire na2190_1;
wire na2191_1;
wire na2192_1;
wire na2193_1;
wire na2194_1;
wire na2195_1;
wire na2196_1;
wire na2197_1;
wire na2198_1;
wire na2199_1;
wire na2200_1;
wire na2201_1;
wire na2202_1;
wire na2203_1;
wire na2204_1;
wire na2205_1;
wire na2206_1;
wire na2207_1;
wire na2208_1;
wire na2209_1;
wire na2210_1;
wire na2211_1;
wire na2212_1;
wire na2213_1;
wire na2214_1;
wire na2215_1;
wire na2216_1;
wire na2217_1;
wire na2218_1;
wire na2219_1;
wire na2220_1;
wire na2221_1;
wire na2222_1;
wire na2223_1;
wire na2224_1;
wire na2225_1;
wire na2226_1;
wire na2227_1;
wire na2228_1;
wire na2229_1;
wire na2230_1;
wire na2231_1;
wire na2232_1;
wire na2233_1;
wire na2234_1;
wire na2235_1;
wire na2236_1;
wire na2237_1;
wire na2238_1;
wire na2239_1;
wire na2240_1;
wire na2241_1;
wire na2242_1;
wire na2243_1;
wire na2244_1;
wire na2245_1;
wire na2246_1;
wire na2247_1;
wire na2248_1;
wire na2249_1;
wire na2250_1;
wire na2251_1;
wire na2252_1;
wire na2253_1;
wire na2254_1;
wire na2255_1;
wire na2256_1;
wire na2257_1;
wire na2258_1;
wire na2259_1;
wire na2260_1;
wire na2261_1;
wire na2262_1;
wire na2263_1;
wire na2264_1;
wire na2265_1;
wire na2266_1;
wire na2267_1;
wire na2268_1;
wire na2269_1;
wire na2270_1;
wire na2271_1;
wire na2272_1;
wire na2273_1;
wire na2274_1;
wire na2275_1;
wire na2276_1;
wire na2277_1;
wire na2278_1;
wire na2279_1;
wire na2280_1;
wire na2281_1;
wire na2282_1;
wire na2283_1;
wire na2284_1;
wire na2285_1;
wire na2286_1;
wire na2287_1;
wire na2288_1;
wire na2289_1;
wire na2290_1;
wire na2291_1;
wire na2292_1;
wire na2293_1;
wire na2294_1;
wire na2295_1;
wire na2296_1;
wire na2297_1;
wire na2298_1;
wire na2299_1;
wire na2300_1;
wire na2301_1;
wire na2302_1;
wire na2303_1;
wire na2304_1;
wire na2305_1;
wire na2306_1;
wire na2307_1;
wire na2308_1;
wire na2309_1;
wire na2310_1;
wire na2311_1;
wire na2312_1;
wire na2313_1;
wire na2314_1;
wire na2315_1;
wire na2316_1;
wire na2317_1;
wire na2318_1;
wire na2319_1;
wire na2320_1;
wire na2321_1;
wire na2322_1;
wire na2323_1;
wire na2324_1;
wire na2325_1;
wire na2326_1;
wire na2327_1;
wire na2328_1;
wire na2329_1;
wire na2330_1;
wire na2331_1;
wire na2332_1;
wire na2333_1;
wire na2334_1;
wire na2335_1;
wire na2336_1;
wire na2337_1;
wire na2338_1;
wire na2339_1;
wire na2340_1;
wire na2341_1;
wire na2342_1;
wire na2343_1;
wire na2344_1;
wire na2345_1;
wire na2346_1;
wire na2347_1;
wire na2348_1;
wire na2349_1;
wire na2350_1;
wire na2351_1;
wire na2352_1;
wire na2353_1;
wire na2354_1;
wire na2355_1;
wire na2356_1;
wire na2357_1;
wire na2358_1;
wire na2359_1;
wire na2360_1;
wire na2361_1;
wire na2362_1;
wire na2363_1;
wire na2364_1;
wire na2365_1;
wire na2366_1;
wire na2367_1;
wire na2368_1;
wire na2369_1;
wire na2370_1;
wire na2371_1;
wire na2372_1;
wire na2373_1;
wire na2374_1;
wire na2375_1;
wire na2376_1;
wire na2377_1;
wire na2378_1;
wire na2379_1;
wire na2380_1;
wire na2381_1;
wire na2382_1;
wire na2383_1;
wire na2384_1;
wire na2385_1;
wire na2386_1;
wire na2387_1;
wire na2388_1;
wire na2389_1;
wire na2390_1;
wire na2401_1;
wire na2402_1;
wire na2403_1;
wire na2404_1;
wire na2405_1;
wire na2406_1;
wire na2407_1;
wire na2408_1;
wire na2409_1;
wire na2410_1;
wire na2411_1;
wire na2412_1;
wire na2412_2;
wire na2413_1;
wire na2414_1;
wire na2415_2;
wire na2416_1;
wire na2417_2;
wire na2422_1;
wire na2422_2;
wire na2423_1;
wire na2425_2;
wire na2426_1;
wire na2431_1;
wire na2431_2;
wire na2432_2;
wire na2434_1;
wire na2435_2;
wire na2440_1;
wire na2440_2;
wire na2441_1;
wire na2443_2;
wire na2444_1;
wire na2449_1;
wire na2449_2;
wire na2450_2;
wire na2452_1;
wire na2453_2;
wire na2458_1;
wire na2458_2;
wire na2459_1;
wire na2461_2;
wire na2462_1;
wire na2467_1;
wire na2467_2;
wire na2468_2;
wire na2470_1;
wire na2471_2;
wire na2476_1;
wire na2476_2;
wire na2477_1;
wire na2479_2;
wire na2480_1;
wire na2485_1;
wire na2485_2;
wire na2486_2;
wire na2488_1;
wire na2489_2;
wire na2494_1;
wire na2494_2;
wire na2495_1;
wire na2497_2;
wire na2498_1;
wire na2503_1;
wire na2504_2;
wire na2505_2;
wire na2506_2;
wire na2507_2;
wire na2508_2;
wire na2509_2;
wire na2510_2;
wire na2511_2;
wire na2512_2;
wire na2513_2;
wire na2514_2;
wire na2515_2;
wire na2516_2;
wire na2517_2;
wire na2518_2;
wire na2519_2;
wire na2520_2;
wire na2521_2;
wire na2522_2;
wire na2523_2;
wire na2524_2;
wire na2504_10;
wire na2505_10;
wire na2506_10;
wire na2507_10;
wire na2508_10;
wire na2509_10;
wire na2510_10;
wire na2511_10;
wire na2512_10;
wire na2513_10;

// C_OR////      x136y42     80'h00_0018_00_0000_0EEE_B7ED
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1_1 ( .OUT(na1_1), .IN1(~na14_1), .IN2(na9_2), .IN3(na2412_1), .IN4(na2416_1), .IN5(~na14_2), .IN6(~na2413_1), .IN7(na2412_2),
                   .IN8(~na2415_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
CLKIN      #(.CLKIN_CFG (32'h0000_0000)) 
           _a2 ( .PCLK0(na2_1), .PCLK1(_d0), .PCLK2(_d1), .PCLK3(_d2), .CLK0(na2390_1), .CLK1(1'b0), .CLK2(1'b0), .CLK3(1'b0), .SER_CLK(1'b0),
                 .SPI_CLK(1'b0), .JTAG_CLK(1'b0) );
// C_AND///AND/      x133y58     80'h00_0078_00_0000_0C88_1244
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4_1 ( .OUT(na4_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2389_1), .IN6(~na2386_1), .IN7(~na2387_1), .IN8(~na2388_1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4_4 ( .OUT(na4_2), .IN1(~na2389_1), .IN2(na2386_1), .IN3(~na2387_1), .IN4(na2388_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                   .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x129y53     80'h00_0078_00_0000_0C88_2441
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5_1 ( .OUT(na5_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2389_1), .IN6(na2386_1), .IN7(na2387_1), .IN8(~na2388_1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5_4 ( .OUT(na5_2), .IN1(~na2389_1), .IN2(~na2386_1), .IN3(~na2387_1), .IN4(na2388_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                   .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x124y57     80'h00_0018_00_0000_0C88_84FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7_1 ( .OUT(na7_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2389_1), .IN6(na2386_1), .IN7(na2387_1), .IN8(na2388_1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x125y46     80'h00_0060_00_0000_0C08_FF5A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9_4 ( .OUT(na9_2), .IN1(na2336_1), .IN2(1'b1), .IN3(~na10_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x124y59     80'h00_0018_00_0040_0CDC_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a10_1 ( .OUT(na10_1), .IN1(1'b1), .IN2(1'b0), .IN3(~na2417_2), .IN4(~na2388_1), .IN5(na2389_1), .IN6(1'b1), .IN7(~na2387_1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x142y53     80'h00_0078_00_0000_0C88_1881
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a12_1 ( .OUT(na12_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2389_1), .IN6(na2386_1), .IN7(~na2387_1), .IN8(~na2388_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a12_4 ( .OUT(na12_2), .IN1(~na2389_1), .IN2(~na2386_1), .IN3(na2387_1), .IN4(na2388_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x139y53     80'h00_0078_00_0000_0C88_2114
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a13_1 ( .OUT(na13_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2389_1), .IN6(~na2386_1), .IN7(na2387_1),
                    .IN8(~na2388_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a13_4 ( .OUT(na13_2), .IN1(~na2389_1), .IN2(na2386_1), .IN3(~na2387_1), .IN4(~na2388_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND///ORAND/      x143y41     80'h00_0078_00_0000_0C88_7777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a14_1 ( .OUT(na14_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na13_2), .IN6(~na1886_1), .IN7(~na12_2), .IN8(~na2136_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a14_4 ( .OUT(na14_2), .IN1(~na13_1), .IN2(~na1936_1), .IN3(~na12_1), .IN4(~na2286_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x137y41     80'h00_0018_00_0000_0EEE_D7DE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a18_1 ( .OUT(na18_1), .IN1(na2426_1), .IN2(na22_1), .IN3(~na24_1), .IN4(na2422_1), .IN5(~na2425_2), .IN6(~na2423_1), .IN7(~na24_2),
                    .IN8(na2422_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x123y46     80'h00_0018_00_0000_0C88_5AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a22_1 ( .OUT(na22_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2341_1), .IN6(1'b1), .IN7(~na10_1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND///ORAND/      x134y47     80'h00_0078_00_0000_0C88_7777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a24_1 ( .OUT(na24_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2091_1), .IN6(~na4_2), .IN7(~na12_1), .IN8(~na2291_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a24_4 ( .OUT(na24_2), .IN1(~na2241_1), .IN2(~na4_1), .IN3(~na12_2), .IN4(~na2141_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x134y48     80'h00_0018_00_0000_0EEE_B7BE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a25_1 ( .OUT(na25_1), .IN1(na2435_2), .IN2(na29_2), .IN3(na2431_1), .IN4(~na31_1), .IN5(~na2434_1), .IN6(~na2432_2), .IN7(na2431_2),
                    .IN8(~na31_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x123y48     80'h00_0060_00_0000_0C08_FF5C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a29_4 ( .OUT(na29_2), .IN1(1'b1), .IN2(na2346_1), .IN3(~na10_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND///ORAND/      x142y48     80'h00_0078_00_0000_0C88_7777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a31_1 ( .OUT(na31_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na13_2), .IN6(~na1896_1), .IN7(~na12_2), .IN8(~na2146_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a31_4 ( .OUT(na31_2), .IN1(~na13_1), .IN2(~na1946_1), .IN3(~na12_1), .IN4(~na2296_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x134y51     80'h00_0018_00_0000_0EEE_D7ED
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a32_1 ( .OUT(na32_1), .IN1(~na38_1), .IN2(na36_1), .IN3(na2444_1), .IN4(na2440_1), .IN5(~na38_2), .IN6(~na2443_2), .IN7(~na2441_1),
                    .IN8(na2440_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x123y50     80'h00_0018_00_0000_0C88_5AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a36_1 ( .OUT(na36_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2351_1), .IN6(1'b1), .IN7(~na10_1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND///ORAND/      x135y53     80'h00_0078_00_0000_0C88_7777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a38_1 ( .OUT(na38_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2101_1), .IN6(~na4_2), .IN7(~na12_1), .IN8(~na2301_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a38_4 ( .OUT(na38_2), .IN1(~na2251_1), .IN2(~na4_1), .IN3(~na12_2), .IN4(~na2151_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x134y53     80'h00_0018_00_0000_0EEE_D7EB
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a39_1 ( .OUT(na39_1), .IN1(na2523_2), .IN2(~na45_1), .IN3(na43_2), .IN4(na2453_2), .IN5(~na2452_1), .IN6(~na45_2), .IN7(~na2450_2),
                    .IN8(na2449_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x124y51     80'h00_0060_00_0000_0C08_FF5C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a43_4 ( .OUT(na43_2), .IN1(1'b1), .IN2(na2356_1), .IN3(~na10_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND///ORAND/      x141y50     80'h00_0078_00_0000_0C88_7777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a45_1 ( .OUT(na45_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na13_2), .IN6(~na1906_1), .IN7(~na12_2), .IN8(~na2156_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a45_4 ( .OUT(na45_2), .IN1(~na13_1), .IN2(~na1956_1), .IN3(~na12_1), .IN4(~na2306_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x137y57     80'h00_0018_00_0000_0EEE_B7BE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a46_1 ( .OUT(na46_1), .IN1(na2462_1), .IN2(na50_1), .IN3(na2458_1), .IN4(~na52_1), .IN5(~na2461_2), .IN6(~na2459_1), .IN7(na2458_2),
                    .IN8(~na52_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x123y60     80'h00_0018_00_0000_0C88_5CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a50_1 ( .OUT(na50_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2361_1), .IN7(~na10_1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND///ORAND/      x142y56     80'h00_0078_00_0000_0C88_7777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a52_1 ( .OUT(na52_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na13_2), .IN6(~na1911_1), .IN7(~na12_2), .IN8(~na2161_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a52_4 ( .OUT(na52_2), .IN1(~na13_1), .IN2(~na1961_1), .IN3(~na12_1), .IN4(~na2311_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x135y63     80'h00_0018_00_0000_0EEE_7DBE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a53_1 ( .OUT(na53_1), .IN1(na57_2), .IN2(na2467_1), .IN3(na2471_2), .IN4(~na59_1), .IN5(~na2468_2), .IN6(na2467_2), .IN7(~na2470_1),
                    .IN8(~na59_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x121y65     80'h00_0060_00_0000_0C08_FF5C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a57_4 ( .OUT(na57_2), .IN1(1'b1), .IN2(na2366_1), .IN3(~na10_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND///ORAND/      x142y58     80'h00_0078_00_0000_0C88_7777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a59_1 ( .OUT(na59_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na13_2), .IN6(~na1916_1), .IN7(~na12_2), .IN8(~na2166_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a59_4 ( .OUT(na59_2), .IN1(~na13_1), .IN2(~na1966_1), .IN3(~na12_1), .IN4(~na2316_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x135y64     80'h00_0018_00_0000_0EEE_B7ED
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a60_1 ( .OUT(na60_1), .IN1(~na66_1), .IN2(na2480_1), .IN3(na2476_1), .IN4(na64_1), .IN5(~na66_2), .IN6(~na2479_2), .IN7(na2476_2),
                    .IN8(~na2477_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x122y66     80'h00_0018_00_0000_0C88_5CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a64_1 ( .OUT(na64_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2371_1), .IN7(~na10_1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND///ORAND/      x145y61     80'h00_0078_00_0000_0C88_7777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a66_1 ( .OUT(na66_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na13_2), .IN6(~na1921_1), .IN7(~na12_2), .IN8(~na2171_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a66_4 ( .OUT(na66_2), .IN1(~na13_1), .IN2(~na1971_1), .IN3(~na12_1), .IN4(~na2321_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x136y66     80'h00_0018_00_0000_0EEE_D7ED
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a67_1 ( .OUT(na67_1), .IN1(~na73_1), .IN2(na71_2), .IN3(na2489_2), .IN4(na2485_1), .IN5(~na73_2), .IN6(~na2488_1), .IN7(~na2486_2),
                    .IN8(na2485_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x125y66     80'h00_0060_00_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a71_4 ( .OUT(na71_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2376_1), .IN4(~na2518_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND///ORAND/      x145y65     80'h00_0078_00_0000_0C88_7777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a73_1 ( .OUT(na73_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na13_2), .IN6(~na1926_1), .IN7(~na12_2), .IN8(~na2176_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a73_4 ( .OUT(na73_2), .IN1(~na13_1), .IN2(~na1976_1), .IN3(~na12_1), .IN4(~na2326_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x136y68     80'h00_0018_00_0000_0EEE_7DED
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a74_1 ( .OUT(na74_1), .IN1(~na80_1), .IN2(na2494_1), .IN3(na78_1), .IN4(na2498_1), .IN5(~na80_2), .IN6(na2494_2), .IN7(~na2495_1),
                    .IN8(~na2497_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x126y67     80'h00_0018_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a78_1 ( .OUT(na78_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2381_1), .IN8(~na2518_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND///ORAND/      x135y65     80'h00_0078_00_0000_0C88_7777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a80_1 ( .OUT(na80_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na5_2), .IN6(~na2081_1), .IN7(~na12_1), .IN8(~na2331_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a80_4 ( .OUT(na80_2), .IN1(~na2281_1), .IN2(~na4_1), .IN3(~na12_2), .IN4(~na2181_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x134y52     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a81_4 ( .OUT(na81_2), .IN1(na82_2), .IN2(1'b1), .IN3(na84_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x131y55     80'h00_0060_00_0000_0C08_FF8C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a82_4 ( .OUT(na82_2), .IN1(1'b1), .IN2(na2521_2), .IN3(na83_1), .IN4(na277_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x134y59     80'h00_0018_00_0000_0C88_48FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a83_1 ( .OUT(na83_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2411_1), .IN6(na2386_1), .IN7(~na2524_2), .IN8(na277_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x128y61     80'h00_0060_00_0000_0C08_FF81
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a84_4 ( .OUT(na84_2), .IN1(~na2384_1), .IN2(~na2383_1), .IN3(na2385_1), .IN4(na2382_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x138y55     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a85_1 ( .OUT(na85_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_2), .IN6(1'b1), .IN7(na86_1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x128y61     80'h00_0018_00_0000_0C88_21FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a86_1 ( .OUT(na86_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2384_1), .IN6(~na2383_1), .IN7(na2385_1),
                    .IN8(~na2382_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x135y49     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a87_4 ( .OUT(na87_2), .IN1(na82_2), .IN2(1'b1), .IN3(na88_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x132y61     80'h00_0018_00_0000_0C88_48FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a88_1 ( .OUT(na88_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2384_1), .IN6(na2383_1), .IN7(~na2385_1), .IN8(na2382_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x141y53     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a89_1 ( .OUT(na89_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_2), .IN6(1'b1), .IN7(na90_1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x128y59     80'h00_0018_00_0000_0C88_42FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a90_1 ( .OUT(na90_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2384_1), .IN6(~na2383_1), .IN7(~na2385_1),
                    .IN8(na2382_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x137y50     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a91_4 ( .OUT(na91_2), .IN1(na82_2), .IN2(1'b1), .IN3(na92_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x130y61     80'h00_0018_00_0000_0C88_18FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a92_1 ( .OUT(na92_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2384_1), .IN6(na2383_1), .IN7(~na2385_1), .IN8(~na2382_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x138y58     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a93_1 ( .OUT(na93_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_2), .IN6(1'b1), .IN7(na94_1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x128y63     80'h00_0018_00_0000_0C88_81FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a94_1 ( .OUT(na94_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2384_1), .IN6(~na2382_1), .IN7(na2385_1),
                    .IN8(na2383_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x135y51     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a95_4 ( .OUT(na95_2), .IN1(na82_2), .IN2(1'b1), .IN3(na96_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x132y57     80'h00_0018_00_0000_0C88_84FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a96_1 ( .OUT(na96_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2384_1), .IN6(na2383_1), .IN7(na2385_1), .IN8(na2382_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x142y54     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a97_1 ( .OUT(na97_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_2), .IN6(1'b1), .IN7(na98_1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x130y59     80'h00_0018_00_0000_0C88_12FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a98_1 ( .OUT(na98_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2384_1), .IN6(~na2383_1), .IN7(~na2385_1),
                    .IN8(~na2382_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x115y64     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a99_4 ( .OUT(na99_2), .IN1(1'b1), .IN2(na100_1), .IN3(na102_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x115y62     80'h00_0018_00_0000_0888_4532
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a100_1 ( .OUT(na100_1), .IN1(na2411_1), .IN2(~na2386_1), .IN3(1'b1), .IN4(~na277_1), .IN5(~na2519_2), .IN6(1'b1), .IN7(~na279_1),
                     .IN8(na2503_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x128y59     80'h00_0060_00_0000_0C08_FF88
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a102_4 ( .OUT(na102_2), .IN1(na2384_1), .IN2(na2383_1), .IN3(na2385_1), .IN4(na2382_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x114y64     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a103_4 ( .OUT(na103_2), .IN1(1'b1), .IN2(na100_1), .IN3(na104_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x126y63     80'h00_0060_00_0000_0C08_FF28
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a104_4 ( .OUT(na104_2), .IN1(na2384_1), .IN2(na2383_1), .IN3(na2385_1), .IN4(~na2382_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x115y63     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a105_4 ( .OUT(na105_2), .IN1(1'b1), .IN2(na100_1), .IN3(na106_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x126y61     80'h00_0060_00_0000_0C08_FF82
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a106_4 ( .OUT(na106_2), .IN1(na2384_1), .IN2(~na2383_1), .IN3(na2385_1), .IN4(na2382_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x140y53     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a107_1 ( .OUT(na107_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_2), .IN6(1'b1), .IN7(na108_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x128y57     80'h00_0060_00_0000_0C08_FF44
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a108_4 ( .OUT(na108_2), .IN1(~na2384_1), .IN2(na2383_1), .IN3(~na2385_1), .IN4(na2382_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x113y63     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a109_4 ( .OUT(na109_2), .IN1(1'b1), .IN2(na100_1), .IN3(na110_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x130y63     80'h00_0018_00_0000_0C88_22FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a110_1 ( .OUT(na110_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2384_1), .IN6(~na2383_1), .IN7(na2385_1),
                     .IN8(~na2382_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x111y62     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a111_1 ( .OUT(na111_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na100_1), .IN7(na96_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x116y66     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a112_4 ( .OUT(na112_2), .IN1(1'b1), .IN2(na100_1), .IN3(na94_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x112y62     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a113_1 ( .OUT(na113_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na100_1), .IN7(na84_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x114y61     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a114_4 ( .OUT(na114_2), .IN1(1'b1), .IN2(na100_1), .IN3(na86_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x138y53     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a115_1 ( .OUT(na115_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_2), .IN6(1'b1), .IN7(na116_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x126y59     80'h00_0018_00_0000_0C88_41FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a116_1 ( .OUT(na116_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2384_1), .IN6(~na2382_1), .IN7(~na2385_1),
                     .IN8(na2383_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x114y58     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a117_4 ( .OUT(na117_2), .IN1(1'b1), .IN2(na100_1), .IN3(na88_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x112y59     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a118_1 ( .OUT(na118_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na100_1), .IN7(na92_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x133y49     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a119_4 ( .OUT(na119_2), .IN1(na82_2), .IN2(1'b1), .IN3(na120_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x126y57     80'h00_0018_00_0000_0C88_41FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a120_1 ( .OUT(na120_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2384_1), .IN6(~na2383_1), .IN7(~na2385_1),
                     .IN8(na2382_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x110y62     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a121_1 ( .OUT(na121_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na100_1), .IN7(na90_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x115y58     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a122_4 ( .OUT(na122_2), .IN1(1'b1), .IN2(na100_1), .IN3(na98_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x142y55     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a123_1 ( .OUT(na123_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_2), .IN6(1'b1), .IN7(na124_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x128y57     80'h00_0018_00_0000_0C88_11FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a124_1 ( .OUT(na124_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2384_1), .IN6(~na2383_1), .IN7(~na2385_1),
                     .IN8(~na2382_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x109y59     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a125_4 ( .OUT(na125_2), .IN1(1'b1), .IN2(na100_1), .IN3(na108_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x110y58     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a126_1 ( .OUT(na126_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na100_1), .IN7(na116_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x113y59     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a127_4 ( .OUT(na127_2), .IN1(1'b1), .IN2(na100_1), .IN3(na120_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x109y58     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a128_1 ( .OUT(na128_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na100_1), .IN7(na124_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x132y55     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a129_4 ( .OUT(na129_2), .IN1(na82_2), .IN2(1'b1), .IN3(na106_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x142y57     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a130_1 ( .OUT(na130_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_2), .IN6(1'b1), .IN7(na110_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x136y53     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a131_4 ( .OUT(na131_2), .IN1(na82_2), .IN2(1'b1), .IN3(na104_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x139y56     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a132_1 ( .OUT(na132_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_2), .IN6(1'b1), .IN7(na102_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x137y47     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a133_4 ( .OUT(na133_2), .IN1(na134_1), .IN2(1'b1), .IN3(na124_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x141y55     80'h00_0018_00_0000_0888_C823
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a134_1 ( .OUT(na134_1), .IN1(1'b1), .IN2(~na2386_1), .IN3(na279_1), .IN4(~na2503_1), .IN5(na2411_1), .IN6(na2520_2), .IN7(1'b1),
                     .IN8(na277_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x141y51     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a136_1 ( .OUT(na136_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na134_1), .IN6(1'b1), .IN7(na120_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x139y52     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a137_4 ( .OUT(na137_2), .IN1(na134_1), .IN2(1'b1), .IN3(na116_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x143y54     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a138_1 ( .OUT(na138_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na134_1), .IN6(1'b1), .IN7(na108_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x137y52     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a139_4 ( .OUT(na139_2), .IN1(na134_1), .IN2(1'b1), .IN3(na98_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x141y58     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a140_1 ( .OUT(na140_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na134_1), .IN6(1'b1), .IN7(na90_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x136y55     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a141_4 ( .OUT(na141_2), .IN1(na134_1), .IN2(1'b1), .IN3(na92_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x145y55     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a142_1 ( .OUT(na142_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na134_1), .IN6(1'b1), .IN7(na88_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x138y54     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a143_4 ( .OUT(na143_2), .IN1(na134_1), .IN2(1'b1), .IN3(na86_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x145y54     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a144_1 ( .OUT(na144_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na134_1), .IN6(1'b1), .IN7(na84_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x140y53     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a145_4 ( .OUT(na145_2), .IN1(na134_1), .IN2(1'b1), .IN3(na94_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x144y54     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a146_1 ( .OUT(na146_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na134_1), .IN6(1'b1), .IN7(na96_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x137y55     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a147_4 ( .OUT(na147_2), .IN1(na134_1), .IN2(1'b1), .IN3(na110_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x145y56     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a148_1 ( .OUT(na148_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na134_1), .IN6(1'b1), .IN7(na106_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x138y56     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a149_4 ( .OUT(na149_2), .IN1(na134_1), .IN2(1'b1), .IN3(na104_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x143y55     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a150_1 ( .OUT(na150_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na134_1), .IN6(1'b1), .IN7(na102_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x120y49     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a151_4 ( .OUT(na151_2), .IN1(na152_1), .IN2(1'b1), .IN3(na124_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x123y53     80'h00_0018_00_0000_0888_382C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a152_1 ( .OUT(na152_1), .IN1(1'b1), .IN2(na2520_2), .IN3(na279_1), .IN4(~na2503_1), .IN5(na2411_1), .IN6(na2386_1), .IN7(1'b1),
                     .IN8(~na277_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x118y52     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a154_1 ( .OUT(na154_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na152_1), .IN6(1'b1), .IN7(na120_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x123y51     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a155_4 ( .OUT(na155_2), .IN1(na152_1), .IN2(1'b1), .IN3(na116_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x121y52     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a156_1 ( .OUT(na156_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na152_1), .IN6(1'b1), .IN7(na108_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x122y50     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a157_4 ( .OUT(na157_2), .IN1(na152_1), .IN2(1'b1), .IN3(na98_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x119y51     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a158_1 ( .OUT(na158_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na152_1), .IN6(1'b1), .IN7(na90_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x123y50     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a159_4 ( .OUT(na159_2), .IN1(na152_1), .IN2(1'b1), .IN3(na92_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x120y52     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a160_1 ( .OUT(na160_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na152_1), .IN6(1'b1), .IN7(na88_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x127y55     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a161_4 ( .OUT(na161_2), .IN1(na152_1), .IN2(1'b1), .IN3(na86_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x123y55     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a162_1 ( .OUT(na162_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na152_1), .IN6(1'b1), .IN7(na84_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x125y58     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a163_4 ( .OUT(na163_2), .IN1(na152_1), .IN2(1'b1), .IN3(na94_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x121y55     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a164_1 ( .OUT(na164_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na152_1), .IN6(1'b1), .IN7(na96_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x124y58     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a165_1 ( .OUT(na165_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na152_1), .IN6(1'b1), .IN7(na110_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x125y55     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a166_1 ( .OUT(na166_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na152_1), .IN6(1'b1), .IN7(na106_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x125y59     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a167_4 ( .OUT(na167_2), .IN1(na152_1), .IN2(1'b1), .IN3(na104_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x122y56     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a168_1 ( .OUT(na168_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na152_1), .IN6(1'b1), .IN7(na102_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x119y57     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a169_4 ( .OUT(na169_2), .IN1(1'b1), .IN2(1'b1), .IN3(na124_1), .IN4(na170_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x128y56     80'h00_0018_00_0000_0888_3A22
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a170_1 ( .OUT(na170_1), .IN1(na2519_2), .IN2(~na2386_1), .IN3(na279_1), .IN4(~na277_1), .IN5(na2411_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(~na2503_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x116y54     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a172_1 ( .OUT(na172_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na120_1), .IN8(na170_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x120y57     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a173_4 ( .OUT(na173_2), .IN1(1'b1), .IN2(1'b1), .IN3(na116_1), .IN4(na170_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x116y55     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a174_1 ( .OUT(na174_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na108_2), .IN8(na170_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x122y58     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a175_4 ( .OUT(na175_2), .IN1(1'b1), .IN2(1'b1), .IN3(na98_1), .IN4(na170_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x118y53     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a176_1 ( .OUT(na176_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na90_1), .IN8(na170_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x123y57     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a177_4 ( .OUT(na177_2), .IN1(1'b1), .IN2(1'b1), .IN3(na92_1), .IN4(na170_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x118y55     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a178_1 ( .OUT(na178_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na88_1), .IN8(na170_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x122y53     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a179_4 ( .OUT(na179_2), .IN1(1'b1), .IN2(1'b1), .IN3(na86_1), .IN4(na170_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x120y54     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a180_1 ( .OUT(na180_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na84_2), .IN8(na170_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x124y53     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a181_4 ( .OUT(na181_2), .IN1(1'b1), .IN2(1'b1), .IN3(na94_1), .IN4(na170_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x119y54     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a182_1 ( .OUT(na182_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na96_1), .IN8(na170_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x121y56     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a183_4 ( .OUT(na183_2), .IN1(1'b1), .IN2(1'b1), .IN3(na110_1), .IN4(na170_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x122y54     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a184_1 ( .OUT(na184_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na106_2), .IN8(na170_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x119y55     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a185_4 ( .OUT(na185_2), .IN1(1'b1), .IN2(1'b1), .IN3(na104_2), .IN4(na170_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x122y53     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a186_1 ( .OUT(na186_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na102_2), .IN8(na170_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x123y61     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a187_4 ( .OUT(na187_2), .IN1(1'b1), .IN2(1'b1), .IN3(na124_1), .IN4(na188_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x128y60     80'h00_0018_00_0000_0C88_2CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a188_1 ( .OUT(na188_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2522_2), .IN7(na83_1), .IN8(~na277_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x127y55     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a189_1 ( .OUT(na189_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na120_1), .IN8(na188_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x125y62     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a190_4 ( .OUT(na190_2), .IN1(1'b1), .IN2(1'b1), .IN3(na116_1), .IN4(na188_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x125y58     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a191_1 ( .OUT(na191_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na108_2), .IN8(na188_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x126y64     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a192_4 ( .OUT(na192_2), .IN1(1'b1), .IN2(1'b1), .IN3(na98_1), .IN4(na188_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x128y55     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a193_1 ( .OUT(na193_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na90_1), .IN8(na188_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x126y59     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a194_4 ( .OUT(na194_2), .IN1(1'b1), .IN2(1'b1), .IN3(na92_1), .IN4(na188_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x126y60     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a195_1 ( .OUT(na195_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na88_1), .IN8(na188_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x123y56     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a196_4 ( .OUT(na196_2), .IN1(1'b1), .IN2(1'b1), .IN3(na86_1), .IN4(na188_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x126y56     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a197_1 ( .OUT(na197_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na84_2), .IN8(na188_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x124y58     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a198_4 ( .OUT(na198_2), .IN1(1'b1), .IN2(1'b1), .IN3(na94_1), .IN4(na188_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x125y54     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a199_1 ( .OUT(na199_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na96_1), .IN8(na188_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x125y61     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a200_4 ( .OUT(na200_2), .IN1(1'b1), .IN2(1'b1), .IN3(na110_1), .IN4(na188_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x128y55     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a201_4 ( .OUT(na201_2), .IN1(1'b1), .IN2(1'b1), .IN3(na106_2), .IN4(na188_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x128y58     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a202_1 ( .OUT(na202_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na104_2), .IN8(na188_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x123y60     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a203_4 ( .OUT(na203_2), .IN1(1'b1), .IN2(1'b1), .IN3(na102_2), .IN4(na188_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x136y60     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a204_4 ( .OUT(na204_2), .IN1(na205_1), .IN2(1'b1), .IN3(na124_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x143y59     80'h00_0018_00_0000_0888_C223
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a205_1 ( .OUT(na205_1), .IN1(1'b1), .IN2(~na2386_1), .IN3(na279_1), .IN4(~na2503_1), .IN5(na2411_1), .IN6(~na2520_2), .IN7(1'b1),
                     .IN8(na277_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x145y59     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a206_1 ( .OUT(na206_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na205_1), .IN6(1'b1), .IN7(na120_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x144y60     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a207_1 ( .OUT(na207_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na205_1), .IN6(1'b1), .IN7(na116_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x145y60     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a208_1 ( .OUT(na208_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na205_1), .IN6(1'b1), .IN7(na108_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x143y58     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a209_1 ( .OUT(na209_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na205_1), .IN6(1'b1), .IN7(na98_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x137y59     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a210_4 ( .OUT(na210_2), .IN1(na205_1), .IN2(1'b1), .IN3(na90_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x146y60     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a211_1 ( .OUT(na211_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na205_1), .IN6(1'b1), .IN7(na92_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x139y59     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a212_4 ( .OUT(na212_2), .IN1(na205_1), .IN2(1'b1), .IN3(na88_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x138y58     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a213_4 ( .OUT(na213_2), .IN1(na205_1), .IN2(1'b1), .IN3(na86_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x146y58     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a214_1 ( .OUT(na214_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na205_1), .IN6(1'b1), .IN7(na84_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x142y57     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a215_4 ( .OUT(na215_2), .IN1(na205_1), .IN2(1'b1), .IN3(na94_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x139y57     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a216_4 ( .OUT(na216_2), .IN1(na205_1), .IN2(1'b1), .IN3(na96_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x138y57     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a217_4 ( .OUT(na217_2), .IN1(na205_1), .IN2(1'b1), .IN3(na110_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x147y60     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a218_1 ( .OUT(na218_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na205_1), .IN6(1'b1), .IN7(na106_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x140y60     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a219_4 ( .OUT(na219_2), .IN1(na205_1), .IN2(1'b1), .IN3(na104_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x145y57     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a220_1 ( .OUT(na220_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na205_1), .IN6(1'b1), .IN7(na102_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x116y60     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a221_4 ( .OUT(na221_2), .IN1(na222_1), .IN2(1'b1), .IN3(na124_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x117y59     80'h00_0018_00_0000_0888_3825
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a222_1 ( .OUT(na222_1), .IN1(~na2519_2), .IN2(1'b1), .IN3(na279_1), .IN4(~na2503_1), .IN5(na2411_1), .IN6(na2386_1), .IN7(1'b1),
                     .IN8(~na277_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x111y57     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a223_1 ( .OUT(na223_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na222_1), .IN6(1'b1), .IN7(na120_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x112y58     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a224_1 ( .OUT(na224_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na222_1), .IN6(1'b1), .IN7(na116_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x116y58     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a225_1 ( .OUT(na225_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na222_1), .IN6(1'b1), .IN7(na108_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x117y60     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a226_4 ( .OUT(na226_2), .IN1(na222_1), .IN2(1'b1), .IN3(na98_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x117y57     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a227_1 ( .OUT(na227_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na222_1), .IN6(1'b1), .IN7(na90_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x119y59     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a228_4 ( .OUT(na228_2), .IN1(na222_1), .IN2(1'b1), .IN3(na92_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x115y58     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a229_1 ( .OUT(na229_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na222_1), .IN6(1'b1), .IN7(na88_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x120y59     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a230_4 ( .OUT(na230_2), .IN1(na222_1), .IN2(1'b1), .IN3(na86_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x114y60     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a231_1 ( .OUT(na231_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na222_1), .IN6(1'b1), .IN7(na84_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x119y61     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a232_4 ( .OUT(na232_2), .IN1(na222_1), .IN2(1'b1), .IN3(na94_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x115y59     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a233_1 ( .OUT(na233_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na222_1), .IN6(1'b1), .IN7(na96_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x118y61     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a234_4 ( .OUT(na234_2), .IN1(na222_1), .IN2(1'b1), .IN3(na110_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x113y60     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a235_1 ( .OUT(na235_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na222_1), .IN6(1'b1), .IN7(na106_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x117y64     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a236_4 ( .OUT(na236_2), .IN1(na222_1), .IN2(1'b1), .IN3(na104_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x116y61     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a237_4 ( .OUT(na237_2), .IN1(na222_1), .IN2(1'b1), .IN3(na102_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x132y60     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a238_4 ( .OUT(na238_2), .IN1(1'b1), .IN2(na239_1), .IN3(na124_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x137y62     80'h00_0018_00_0000_0888_3223
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a239_1 ( .OUT(na239_1), .IN1(1'b1), .IN2(~na2386_1), .IN3(na279_1), .IN4(~na277_1), .IN5(na2411_1), .IN6(~na2520_2), .IN7(1'b1),
                     .IN8(~na2503_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x135y57     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a240_1 ( .OUT(na240_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na239_1), .IN7(na120_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x130y59     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a241_4 ( .OUT(na241_2), .IN1(1'b1), .IN2(na239_1), .IN3(na116_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x135y58     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a242_1 ( .OUT(na242_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na239_1), .IN7(na108_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x127y59     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a243_4 ( .OUT(na243_2), .IN1(1'b1), .IN2(na239_1), .IN3(na98_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x132y59     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a244_1 ( .OUT(na244_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na239_1), .IN7(na90_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x129y59     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a245_4 ( .OUT(na245_2), .IN1(1'b1), .IN2(na239_1), .IN3(na92_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x133y61     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a246_1 ( .OUT(na246_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na239_1), .IN7(na88_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x131y57     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a247_4 ( .OUT(na247_2), .IN1(1'b1), .IN2(na239_1), .IN3(na86_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x135y62     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a248_1 ( .OUT(na248_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na239_1), .IN7(na84_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x131y60     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a249_4 ( .OUT(na249_2), .IN1(1'b1), .IN2(na239_1), .IN3(na94_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x134y62     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a250_1 ( .OUT(na250_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na239_1), .IN7(na96_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x133y60     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a251_1 ( .OUT(na251_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na239_1), .IN7(na110_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x137y60     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a252_1 ( .OUT(na252_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na239_1), .IN7(na106_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x132y58     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a253_4 ( .OUT(na253_2), .IN1(1'b1), .IN2(na239_1), .IN3(na104_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x133y57     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a254_1 ( .OUT(na254_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na239_1), .IN7(na102_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x139y56     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a255_4 ( .OUT(na255_2), .IN1(1'b1), .IN2(1'b1), .IN3(na124_1), .IN4(na256_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x144y58     80'h00_0018_00_0000_0C88_83FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a256_1 ( .OUT(na256_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na2521_2), .IN7(na83_1), .IN8(na277_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x146y56     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a257_1 ( .OUT(na257_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na120_1), .IN8(na256_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x142y55     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a258_4 ( .OUT(na258_2), .IN1(1'b1), .IN2(1'b1), .IN3(na116_1), .IN4(na256_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x147y56     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a259_1 ( .OUT(na259_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na108_2), .IN8(na256_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x138y61     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a260_4 ( .OUT(na260_2), .IN1(1'b1), .IN2(1'b1), .IN3(na98_1), .IN4(na256_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x150y55     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a261_1 ( .OUT(na261_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na90_1), .IN8(na256_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x143y61     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a262_4 ( .OUT(na262_2), .IN1(1'b1), .IN2(1'b1), .IN3(na92_1), .IN4(na256_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x149y56     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a263_1 ( .OUT(na263_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na88_1), .IN8(na256_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x142y54     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a264_4 ( .OUT(na264_2), .IN1(1'b1), .IN2(1'b1), .IN3(na86_1), .IN4(na256_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x141y64     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a265_4 ( .OUT(na265_2), .IN1(1'b1), .IN2(1'b1), .IN3(na84_2), .IN4(na256_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x141y60     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a266_4 ( .OUT(na266_2), .IN1(1'b1), .IN2(1'b1), .IN3(na94_1), .IN4(na256_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x148y56     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a267_1 ( .OUT(na267_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na96_1), .IN8(na256_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x145y63     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a268_4 ( .OUT(na268_2), .IN1(1'b1), .IN2(1'b1), .IN3(na110_1), .IN4(na256_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x147y58     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a269_1 ( .OUT(na269_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na106_2), .IN8(na256_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x144y64     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a270_4 ( .OUT(na270_2), .IN1(1'b1), .IN2(1'b1), .IN3(na104_2), .IN4(na256_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x150y56     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a271_1 ( .OUT(na271_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na102_2), .IN8(na256_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x130y56     80'h00_0078_00_0020_0C66_5330
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a277_1 ( .OUT(na277_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na2386_1), .IN7(~na2387_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na280_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a277_4 ( .OUT(na277_2), .COUTY1(na277_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na2388_1), .IN5(1'b1), .IN6(~na2386_1),
                     .IN7(~na2387_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na280_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x130y57     80'h00_0018_00_0010_0666_0005
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a279_1 ( .OUT(na279_1), .COUTY1(na279_4), .IN1(~na2389_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na277_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x130y55     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a280_2 ( .OUT(na280_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a280_6 ( .COUTY1(na280_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na280_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/D      x136y32     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a282_4 ( .OUT(na282_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a282_5 ( .OUT(na282_2), .CLK(na2414_1), .EN(na97_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na282_2_i) );
// C_AND/D///      x137y31     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a283_1 ( .OUT(na283_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a283_2 ( .OUT(na283_1), .CLK(na2414_1), .EN(na97_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na283_1_i) );
// C_AND/D///      x146y40     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a284_1 ( .OUT(na284_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2403_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a284_2 ( .OUT(na284_1), .CLK(na2414_1), .EN(na97_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na284_1_i) );
// C_AND/D///      x127y46     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a285_1 ( .OUT(na285_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a285_2 ( .OUT(na285_1), .CLK(na2414_1), .EN(na97_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na285_1_i) );
// C_///AND/D      x136y49     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a286_4 ( .OUT(na286_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a286_5 ( .OUT(na286_2), .CLK(na2414_1), .EN(na97_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na286_2_i) );
// C_///AND/D      x142y49     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a287_4 ( .OUT(na287_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2406_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a287_5 ( .OUT(na287_2), .CLK(na2414_1), .EN(na97_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na287_2_i) );
// C_///AND/D      x130y60     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a288_4 ( .OUT(na288_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a288_5 ( .OUT(na288_2), .CLK(na2414_1), .EN(na97_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na288_2_i) );
// C_AND/D///      x142y67     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a289_1 ( .OUT(na289_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a289_2 ( .OUT(na289_1), .CLK(na2414_1), .EN(na97_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na289_1_i) );
// C_AND/D///      x142y73     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a290_1 ( .OUT(na290_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2409_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a290_2 ( .OUT(na290_1), .CLK(na2414_1), .EN(na97_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na290_1_i) );
// C_AND/D///      x133y75     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a291_1 ( .OUT(na291_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a291_2 ( .OUT(na291_1), .CLK(na2414_1), .EN(na97_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na291_1_i) );
// C_///AND/D      x142y35     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a292_4 ( .OUT(na292_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a292_5 ( .OUT(na292_2), .CLK(na2414_1), .EN(na131_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na292_2_i) );
// C_AND/D///      x146y33     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a293_1 ( .OUT(na293_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a293_2 ( .OUT(na293_1), .CLK(na2414_1), .EN(na131_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na293_1_i) );
// C_///AND/D      x139y41     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a294_4 ( .OUT(na294_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a294_5 ( .OUT(na294_2), .CLK(na2414_1), .EN(na131_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na294_2_i) );
// C_///AND/D      x124y47     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a295_4 ( .OUT(na295_2_i), .IN1(1'b1), .IN2(na2404_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a295_5 ( .OUT(na295_2), .CLK(na2414_1), .EN(na131_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na295_2_i) );
// C_///AND/D      x146y57     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a296_4 ( .OUT(na296_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a296_5 ( .OUT(na296_2), .CLK(na2414_1), .EN(na131_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na296_2_i) );
// C_AND/D///      x148y53     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a297_1 ( .OUT(na297_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a297_2 ( .OUT(na297_1), .CLK(na2414_1), .EN(na131_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na297_1_i) );
// C_AND/D///      x140y61     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a298_1 ( .OUT(na298_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2407_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a298_2 ( .OUT(na298_1), .CLK(na2414_1), .EN(na131_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na298_1_i) );
// C_AND/D///      x139y67     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a299_1 ( .OUT(na299_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a299_2 ( .OUT(na299_1), .CLK(na2414_1), .EN(na131_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na299_1_i) );
// C_///AND/D      x142y79     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a300_4 ( .OUT(na300_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a300_5 ( .OUT(na300_2), .CLK(na2414_1), .EN(na131_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na300_2_i) );
// C_///AND/D      x134y84     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a301_4 ( .OUT(na301_2_i), .IN1(1'b1), .IN2(na2410_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a301_5 ( .OUT(na301_2), .CLK(na2414_1), .EN(na131_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na301_2_i) );
// C_///AND/D      x139y34     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a302_4 ( .OUT(na302_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a302_5 ( .OUT(na302_2), .CLK(na2414_1), .EN(na129_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na302_2_i) );
// C_AND/D///      x147y34     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a303_1 ( .OUT(na303_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a303_2 ( .OUT(na303_1), .CLK(na2414_1), .EN(na129_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na303_1_i) );
// C_///AND/D      x136y44     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a304_4 ( .OUT(na304_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a304_5 ( .OUT(na304_2), .CLK(na2414_1), .EN(na129_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na304_2_i) );
// C_AND/D///      x123y48     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a305_1 ( .OUT(na305_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a305_2 ( .OUT(na305_1), .CLK(na2414_1), .EN(na129_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na305_1_i) );
// C_AND/D///      x151y48     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a306_1 ( .OUT(na306_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2405_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a306_2 ( .OUT(na306_1), .CLK(na2414_1), .EN(na129_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na306_1_i) );
// C_AND/D///      x149y54     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a307_1 ( .OUT(na307_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a307_2 ( .OUT(na307_1), .CLK(na2414_1), .EN(na129_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na307_1_i) );
// C_///AND/D      x133y62     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a308_4 ( .OUT(na308_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a308_5 ( .OUT(na308_2), .CLK(na2414_1), .EN(na129_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na308_2_i) );
// C_///AND/D      x142y72     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a309_4 ( .OUT(na309_2_i), .IN1(na2408_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a309_5 ( .OUT(na309_2), .CLK(na2414_1), .EN(na129_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na309_2_i) );
// C_///AND/D      x143y80     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a310_4 ( .OUT(na310_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a310_5 ( .OUT(na310_2), .CLK(na2414_1), .EN(na129_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na310_2_i) );
// C_AND/D///      x135y77     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a311_1 ( .OUT(na311_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a311_2 ( .OUT(na311_1), .CLK(na2414_1), .EN(na129_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na311_1_i) );
// C_AND/D///      x147y37     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a312_1 ( .OUT(na312_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2401_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a312_2 ( .OUT(na312_1), .CLK(na2414_1), .EN(na130_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na312_1_i) );
// C_AND/D///      x147y39     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a313_1 ( .OUT(na313_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a313_2 ( .OUT(na313_1), .CLK(na2414_1), .EN(na130_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na313_1_i) );
// C_///AND/D      x136y41     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a314_4 ( .OUT(na314_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a314_5 ( .OUT(na314_2), .CLK(na2414_1), .EN(na130_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na314_2_i) );
// C_AND/D///      x125y47     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a315_1 ( .OUT(na315_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a315_2 ( .OUT(na315_1), .CLK(na2414_1), .EN(na130_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na315_1_i) );
// C_///AND/D      x147y57     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a316_4 ( .OUT(na316_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a316_5 ( .OUT(na316_2), .CLK(na2414_1), .EN(na130_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na316_2_i) );
// C_///AND/D      x145y59     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a317_4 ( .OUT(na317_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2406_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a317_5 ( .OUT(na317_2), .CLK(na2414_1), .EN(na130_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na317_2_i) );
// C_///AND/D      x137y61     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a318_4 ( .OUT(na318_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a318_5 ( .OUT(na318_2), .CLK(na2414_1), .EN(na130_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na318_2_i) );
// C_AND/D///      x140y67     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a319_1 ( .OUT(na319_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a319_2 ( .OUT(na319_1), .CLK(na2414_1), .EN(na130_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na319_1_i) );
// C_AND/D///      x145y75     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a320_1 ( .OUT(na320_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2409_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a320_2 ( .OUT(na320_1), .CLK(na2414_1), .EN(na130_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na320_1_i) );
// C_AND/D///      x135y78     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a321_1 ( .OUT(na321_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a321_2 ( .OUT(na321_1), .CLK(na2414_1), .EN(na130_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na321_1_i) );
// C_///AND/D      x141y38     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a322_4 ( .OUT(na322_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a322_5 ( .OUT(na322_2), .CLK(na2414_1), .EN(na95_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na322_2_i) );
// C_///AND/D      x136y36     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a323_4 ( .OUT(na323_2_i), .IN1(na2402_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a323_5 ( .OUT(na323_2), .CLK(na2414_1), .EN(na95_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na323_2_i) );
// C_///AND/D      x136y39     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a324_4 ( .OUT(na324_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a324_5 ( .OUT(na324_2), .CLK(na2414_1), .EN(na95_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na324_2_i) );
// C_AND/D///      x121y46     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a325_1 ( .OUT(na325_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a325_2 ( .OUT(na325_1), .CLK(na2414_1), .EN(na95_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na325_1_i) );
// C_///AND/D      x144y57     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a326_4 ( .OUT(na326_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a326_5 ( .OUT(na326_2), .CLK(na2414_1), .EN(na95_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na326_2_i) );
// C_AND/D///      x145y50     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a327_1 ( .OUT(na327_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a327_2 ( .OUT(na327_1), .CLK(na2414_1), .EN(na95_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na327_1_i) );
// C_AND/D///      x141y64     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a328_1 ( .OUT(na328_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2407_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a328_2 ( .OUT(na328_1), .CLK(na2414_1), .EN(na95_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na328_1_i) );
// C_AND/D///      x139y66     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a329_1 ( .OUT(na329_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a329_2 ( .OUT(na329_1), .CLK(na2414_1), .EN(na95_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na329_1_i) );
// C_///AND/D      x136y73     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a330_4 ( .OUT(na330_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a330_5 ( .OUT(na330_2), .CLK(na2414_1), .EN(na95_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na330_2_i) );
// C_///AND/D      x128y82     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a331_4 ( .OUT(na331_2_i), .IN1(1'b1), .IN2(na2410_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a331_5 ( .OUT(na331_2), .CLK(na2414_1), .EN(na95_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na331_2_i) );
// C_///AND/D      x139y39     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a332_4 ( .OUT(na332_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a332_5 ( .OUT(na332_2), .CLK(na2414_1), .EN(na93_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na332_2_i) );
// C_AND/D///      x136y31     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a333_1 ( .OUT(na333_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a333_2 ( .OUT(na333_1), .CLK(na2414_1), .EN(na93_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na333_1_i) );
// C_AND/D///      x144y40     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a334_1 ( .OUT(na334_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2403_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a334_2 ( .OUT(na334_1), .CLK(na2414_1), .EN(na93_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na334_1_i) );
// C_AND/D///      x121y47     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a335_1 ( .OUT(na335_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a335_2 ( .OUT(na335_1), .CLK(na2414_1), .EN(na93_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na335_1_i) );
// C_///AND/D      x146y58     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a336_4 ( .OUT(na336_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a336_5 ( .OUT(na336_2), .CLK(na2414_1), .EN(na93_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na336_2_i) );
// C_AND/D///      x145y49     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a337_1 ( .OUT(na337_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a337_2 ( .OUT(na337_1), .CLK(na2414_1), .EN(na93_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na337_1_i) );
// C_///AND/D      x139y61     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a338_4 ( .OUT(na338_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a338_5 ( .OUT(na338_2), .CLK(na2414_1), .EN(na93_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na338_2_i) );
// C_///AND/D      x139y69     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a339_4 ( .OUT(na339_2_i), .IN1(na2408_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a339_5 ( .OUT(na339_2), .CLK(na2414_1), .EN(na93_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na339_2_i) );
// C_///AND/D      x142y74     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a340_4 ( .OUT(na340_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a340_5 ( .OUT(na340_2), .CLK(na2414_1), .EN(na93_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na340_2_i) );
// C_AND/D///      x122y81     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a341_1 ( .OUT(na341_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a341_2 ( .OUT(na341_1), .CLK(na2414_1), .EN(na93_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na341_1_i) );
// C_AND/D///      x148y33     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a342_1 ( .OUT(na342_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2401_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a342_2 ( .OUT(na342_1), .CLK(na2414_1), .EN(na89_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na342_1_i) );
// C_AND/D///      x141y32     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a343_1 ( .OUT(na343_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a343_2 ( .OUT(na343_1), .CLK(na2414_1), .EN(na89_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na343_1_i) );
// C_///AND/D      x138y39     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a344_4 ( .OUT(na344_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a344_5 ( .OUT(na344_2), .CLK(na2414_1), .EN(na89_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na344_2_i) );
// C_///AND/D      x127y45     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a345_4 ( .OUT(na345_2_i), .IN1(1'b1), .IN2(na2404_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a345_5 ( .OUT(na345_2), .CLK(na2414_1), .EN(na89_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na345_2_i) );
// C_///AND/D      x136y50     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a346_4 ( .OUT(na346_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a346_5 ( .OUT(na346_2), .CLK(na2414_1), .EN(na89_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na346_2_i) );
// C_AND/D///      x144y48     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a347_1 ( .OUT(na347_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a347_2 ( .OUT(na347_1), .CLK(na2414_1), .EN(na89_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na347_1_i) );
// C_///AND/D      x134y59     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a348_4 ( .OUT(na348_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a348_5 ( .OUT(na348_2), .CLK(na2414_1), .EN(na89_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na348_2_i) );
// C_AND/D///      x146y66     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a349_1 ( .OUT(na349_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a349_2 ( .OUT(na349_1), .CLK(na2414_1), .EN(na89_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na349_1_i) );
// C_AND/D///      x144y74     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a350_1 ( .OUT(na350_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2409_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a350_2 ( .OUT(na350_1), .CLK(na2414_1), .EN(na89_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na350_1_i) );
// C_AND/D///      x131y78     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a351_1 ( .OUT(na351_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a351_2 ( .OUT(na351_1), .CLK(na2414_1), .EN(na89_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na351_1_i) );
// C_///AND/D      x136y30     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a352_4 ( .OUT(na352_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a352_5 ( .OUT(na352_2), .CLK(na2414_1), .EN(na107_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na352_2_i) );
// C_///AND/D      x136y37     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a353_4 ( .OUT(na353_2_i), .IN1(na2402_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a353_5 ( .OUT(na353_2), .CLK(na2414_1), .EN(na107_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na353_2_i) );
// C_///AND/D      x139y37     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a354_4 ( .OUT(na354_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a354_5 ( .OUT(na354_2), .CLK(na2414_1), .EN(na107_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na354_2_i) );
// C_AND/D///      x124y46     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a355_1 ( .OUT(na355_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a355_2 ( .OUT(na355_1), .CLK(na2414_1), .EN(na107_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na355_1_i) );
// C_AND/D///      x148y46     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a356_1 ( .OUT(na356_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2405_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a356_2 ( .OUT(na356_1), .CLK(na2414_1), .EN(na107_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na356_1_i) );
// C_AND/D///      x144y52     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a357_1 ( .OUT(na357_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a357_2 ( .OUT(na357_1), .CLK(na2414_1), .EN(na107_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na357_1_i) );
// C_///AND/D      x135y58     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a358_4 ( .OUT(na358_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a358_5 ( .OUT(na358_2), .CLK(na2414_1), .EN(na107_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na358_2_i) );
// C_AND/D///      x143y68     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a359_1 ( .OUT(na359_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a359_2 ( .OUT(na359_1), .CLK(na2414_1), .EN(na107_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na359_1_i) );
// C_///AND/D      x143y78     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a360_4 ( .OUT(na360_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a360_5 ( .OUT(na360_2), .CLK(na2414_1), .EN(na107_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na360_2_i) );
// C_///AND/D      x132y84     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a361_4 ( .OUT(na361_2_i), .IN1(1'b1), .IN2(na2410_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a361_5 ( .OUT(na361_2), .CLK(na2414_1), .EN(na107_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na361_2_i) );
// C_///AND/D      x137y35     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a362_4 ( .OUT(na362_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a362_5 ( .OUT(na362_2), .CLK(na2414_1), .EN(na123_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na362_2_i) );
// C_AND/D///      x141y36     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a363_1 ( .OUT(na363_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a363_2 ( .OUT(na363_1), .CLK(na2414_1), .EN(na123_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na363_1_i) );
// C_AND/D///      x146y38     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a364_1 ( .OUT(na364_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2403_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a364_2 ( .OUT(na364_1), .CLK(na2414_1), .EN(na123_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na364_1_i) );
// C_AND/D///      x125y43     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a365_1 ( .OUT(na365_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a365_2 ( .OUT(na365_1), .CLK(na2414_1), .EN(na123_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na365_1_i) );
// C_///AND/D      x139y45     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a366_4 ( .OUT(na366_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a366_5 ( .OUT(na366_2), .CLK(na2414_1), .EN(na123_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na366_2_i) );
// C_///AND/D      x141y51     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a367_4 ( .OUT(na367_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2406_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a367_5 ( .OUT(na367_2), .CLK(na2414_1), .EN(na123_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na367_2_i) );
// C_///AND/D      x136y57     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a368_4 ( .OUT(na368_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a368_5 ( .OUT(na368_2), .CLK(na2414_1), .EN(na123_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na368_2_i) );
// C_AND/D///      x144y65     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a369_1 ( .OUT(na369_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a369_2 ( .OUT(na369_1), .CLK(na2414_1), .EN(na123_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na369_1_i) );
// C_///AND/D      x148y77     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a370_4 ( .OUT(na370_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a370_5 ( .OUT(na370_2), .CLK(na2414_1), .EN(na123_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na370_2_i) );
// C_AND/D///      x133y81     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a371_1 ( .OUT(na371_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a371_2 ( .OUT(na371_1), .CLK(na2414_1), .EN(na123_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na371_1_i) );
// C_AND/D///      x150y37     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a372_1 ( .OUT(na372_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2401_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a372_2 ( .OUT(na372_1), .CLK(na2414_1), .EN(na85_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na372_1_i) );
// C_AND/D///      x135y31     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a373_1 ( .OUT(na373_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a373_2 ( .OUT(na373_1), .CLK(na2414_1), .EN(na85_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na373_1_i) );
// C_///AND/D      x133y42     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a374_4 ( .OUT(na374_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a374_5 ( .OUT(na374_2), .CLK(na2414_1), .EN(na85_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na374_2_i) );
// C_///AND/D      x124y45     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a375_4 ( .OUT(na375_2_i), .IN1(1'b1), .IN2(na2404_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a375_5 ( .OUT(na375_2), .CLK(na2414_1), .EN(na85_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na375_2_i) );
// C_///AND/D      x143y58     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a376_4 ( .OUT(na376_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a376_5 ( .OUT(na376_2), .CLK(na2414_1), .EN(na85_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na376_2_i) );
// C_AND/D///      x146y51     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a377_1 ( .OUT(na377_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a377_2 ( .OUT(na377_1), .CLK(na2414_1), .EN(na85_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na377_1_i) );
// C_AND/D///      x142y63     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a378_1 ( .OUT(na378_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2407_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a378_2 ( .OUT(na378_1), .CLK(na2414_1), .EN(na85_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na378_1_i) );
// C_AND/D///      x140y65     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a379_1 ( .OUT(na379_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a379_2 ( .OUT(na379_1), .CLK(na2414_1), .EN(na85_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na379_1_i) );
// C_///AND/D      x139y74     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a380_4 ( .OUT(na380_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a380_5 ( .OUT(na380_2), .CLK(na2414_1), .EN(na85_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na380_2_i) );
// C_AND/D///      x123y81     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a381_1 ( .OUT(na381_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a381_2 ( .OUT(na381_1), .CLK(na2414_1), .EN(na85_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na381_1_i) );
// C_///AND/D      x139y33     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a382_4 ( .OUT(na382_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a382_5 ( .OUT(na382_2), .CLK(na2414_1), .EN(na87_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na382_2_i) );
// C_///AND/D      x134y34     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a383_4 ( .OUT(na383_2_i), .IN1(na2402_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a383_5 ( .OUT(na383_2), .CLK(na2414_1), .EN(na87_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na383_2_i) );
// C_///AND/D      x139y43     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a384_4 ( .OUT(na384_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a384_5 ( .OUT(na384_2), .CLK(na2414_1), .EN(na87_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na384_2_i) );
// C_AND/D///      x130y47     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a385_1 ( .OUT(na385_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a385_2 ( .OUT(na385_1), .CLK(na2414_1), .EN(na87_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na385_1_i) );
// C_AND/D///      x145y48     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a386_1 ( .OUT(na386_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2405_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a386_2 ( .OUT(na386_1), .CLK(na2414_1), .EN(na87_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na386_1_i) );
// C_AND/D///      x141y52     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a387_1 ( .OUT(na387_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a387_2 ( .OUT(na387_1), .CLK(na2414_1), .EN(na87_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na387_1_i) );
// C_///AND/D      x133y59     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a388_4 ( .OUT(na388_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a388_5 ( .OUT(na388_2), .CLK(na2414_1), .EN(na87_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na388_2_i) );
// C_///AND/D      x141y70     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a389_4 ( .OUT(na389_2_i), .IN1(na2408_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a389_5 ( .OUT(na389_2), .CLK(na2414_1), .EN(na87_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na389_2_i) );
// C_///AND/D      x141y76     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a390_4 ( .OUT(na390_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a390_5 ( .OUT(na390_2), .CLK(na2414_1), .EN(na87_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na390_2_i) );
// C_AND/D///      x132y80     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a391_1 ( .OUT(na391_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a391_2 ( .OUT(na391_1), .CLK(na2414_1), .EN(na87_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na391_1_i) );
// C_///AND/D      x141y34     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a392_4 ( .OUT(na392_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a392_5 ( .OUT(na392_2), .CLK(na2414_1), .EN(na91_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na392_2_i) );
// C_AND/D///      x142y31     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a393_1 ( .OUT(na393_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a393_2 ( .OUT(na393_1), .CLK(na2414_1), .EN(na91_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na393_1_i) );
// C_AND/D///      x147y40     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a394_1 ( .OUT(na394_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2403_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a394_2 ( .OUT(na394_1), .CLK(na2414_1), .EN(na91_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na394_1_i) );
// C_AND/D///      x130y48     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a395_1 ( .OUT(na395_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a395_2 ( .OUT(na395_1), .CLK(na2414_1), .EN(na91_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na395_1_i) );
// C_///AND/D      x139y47     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a396_4 ( .OUT(na396_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a396_5 ( .OUT(na396_2), .CLK(na2414_1), .EN(na91_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na396_2_i) );
// C_///AND/D      x139y49     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a397_4 ( .OUT(na397_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2406_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a397_5 ( .OUT(na397_2), .CLK(na2414_1), .EN(na91_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na397_2_i) );
// C_///AND/D      x137y60     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a398_4 ( .OUT(na398_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a398_5 ( .OUT(na398_2), .CLK(na2414_1), .EN(na91_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na398_2_i) );
// C_AND/D///      x145y67     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a399_1 ( .OUT(na399_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a399_2 ( .OUT(na399_1), .CLK(na2414_1), .EN(na91_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na399_1_i) );
// C_AND/D///      x143y75     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a400_1 ( .OUT(na400_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2409_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a400_2 ( .OUT(na400_1), .CLK(na2414_1), .EN(na91_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na400_1_i) );
// C_AND/D///      x136y77     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a401_1 ( .OUT(na401_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a401_2 ( .OUT(na401_1), .CLK(na2414_1), .EN(na91_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na401_1_i) );
// C_///AND/D      x106y34     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a402_4 ( .OUT(na402_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a402_5 ( .OUT(na402_2), .CLK(na2414_1), .EN(na128_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na402_2_i) );
// C_AND/D///      x105y37     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a403_1 ( .OUT(na403_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a403_2 ( .OUT(na403_1), .CLK(na2414_1), .EN(na128_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na403_1_i) );
// C_///AND/D      x109y45     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a404_4 ( .OUT(na404_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a404_5 ( .OUT(na404_2), .CLK(na2414_1), .EN(na128_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na404_2_i) );
// C_///AND/D      x113y49     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a405_4 ( .OUT(na405_2_i), .IN1(1'b1), .IN2(na2404_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a405_5 ( .OUT(na405_2), .CLK(na2414_1), .EN(na128_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na405_2_i) );
// C_///AND/D      x107y53     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a406_4 ( .OUT(na406_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a406_5 ( .OUT(na406_2), .CLK(na2414_1), .EN(na128_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na406_2_i) );
// C_AND/D///      x106y61     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a407_1 ( .OUT(na407_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a407_2 ( .OUT(na407_1), .CLK(na2414_1), .EN(na128_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na407_1_i) );
// C_AND/D///      x105y70     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a408_1 ( .OUT(na408_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2407_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a408_2 ( .OUT(na408_1), .CLK(na2414_1), .EN(na128_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na408_1_i) );
// C_AND/D///      x107y77     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a409_1 ( .OUT(na409_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a409_2 ( .OUT(na409_1), .CLK(na2414_1), .EN(na128_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na409_1_i) );
// C_///AND/D      x111y73     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a410_4 ( .OUT(na410_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a410_5 ( .OUT(na410_2), .CLK(na2414_1), .EN(na128_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na410_2_i) );
// C_///AND/D      x127y81     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a411_4 ( .OUT(na411_2_i), .IN1(1'b1), .IN2(na2410_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a411_5 ( .OUT(na411_2), .CLK(na2414_1), .EN(na128_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na411_2_i) );
// C_///AND/D      x138y35     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a412_4 ( .OUT(na412_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a412_5 ( .OUT(na412_2), .CLK(na2414_1), .EN(na115_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na412_2_i) );
// C_AND/D///      x142y34     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a413_1 ( .OUT(na413_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a413_2 ( .OUT(na413_1), .CLK(na2414_1), .EN(na115_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na413_1_i) );
// C_///AND/D      x137y38     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a414_4 ( .OUT(na414_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a414_5 ( .OUT(na414_2), .CLK(na2414_1), .EN(na115_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na414_2_i) );
// C_AND/D///      x128y45     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a415_1 ( .OUT(na415_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a415_2 ( .OUT(na415_1), .CLK(na2414_1), .EN(na115_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na415_1_i) );
// C_AND/D///      x148y45     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a416_1 ( .OUT(na416_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2405_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a416_2 ( .OUT(na416_1), .CLK(na2414_1), .EN(na115_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na416_1_i) );
// C_AND/D///      x146y53     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a417_1 ( .OUT(na417_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a417_2 ( .OUT(na417_1), .CLK(na2414_1), .EN(na115_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na417_1_i) );
// C_///AND/D      x133y57     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a418_4 ( .OUT(na418_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a418_5 ( .OUT(na418_2), .CLK(na2414_1), .EN(na115_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na418_2_i) );
// C_///AND/D      x139y71     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a419_4 ( .OUT(na419_2_i), .IN1(na2408_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a419_5 ( .OUT(na419_2), .CLK(na2414_1), .EN(na115_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na419_2_i) );
// C_///AND/D      x139y77     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a420_4 ( .OUT(na420_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a420_5 ( .OUT(na420_2), .CLK(na2414_1), .EN(na115_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na420_2_i) );
// C_AND/D///      x130y81     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a421_1 ( .OUT(na421_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a421_2 ( .OUT(na421_1), .CLK(na2414_1), .EN(na115_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na421_1_i) );
// C_AND/D///      x143y36     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a422_1 ( .OUT(na422_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2401_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a422_2 ( .OUT(na422_1), .CLK(na2414_1), .EN(na119_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na422_1_i) );
// C_AND/D///      x143y33     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a423_1 ( .OUT(na423_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a423_2 ( .OUT(na423_1), .CLK(na2414_1), .EN(na119_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na423_1_i) );
// C_///AND/D      x138y37     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a424_4 ( .OUT(na424_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a424_5 ( .OUT(na424_2), .CLK(na2414_1), .EN(na119_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na424_2_i) );
// C_AND/D///      x129y46     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a425_1 ( .OUT(na425_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a425_2 ( .OUT(na425_1), .CLK(na2414_1), .EN(na119_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na425_1_i) );
// C_///AND/D      x141y48     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a426_4 ( .OUT(na426_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a426_5 ( .OUT(na426_2), .CLK(na2414_1), .EN(na119_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na426_2_i) );
// C_///AND/D      x139y54     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a427_4 ( .OUT(na427_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2406_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a427_5 ( .OUT(na427_2), .CLK(na2414_1), .EN(na119_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na427_2_i) );
// C_///AND/D      x136y58     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a428_4 ( .OUT(na428_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a428_5 ( .OUT(na428_2), .CLK(na2414_1), .EN(na119_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na428_2_i) );
// C_AND/D///      x142y70     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a429_1 ( .OUT(na429_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a429_2 ( .OUT(na429_1), .CLK(na2414_1), .EN(na119_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na429_1_i) );
// C_AND/D///      x146y76     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a430_1 ( .OUT(na430_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2409_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a430_2 ( .OUT(na430_1), .CLK(na2414_1), .EN(na119_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na430_1_i) );
// C_AND/D///      x131y82     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a431_1 ( .OUT(na431_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a431_2 ( .OUT(na431_1), .CLK(na2414_1), .EN(na119_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na431_1_i) );
// C_///AND/D      x144y38     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a432_4 ( .OUT(na432_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a432_5 ( .OUT(na432_2), .CLK(na2414_1), .EN(na132_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na432_2_i) );
// C_///AND/D      x138y42     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a433_4 ( .OUT(na433_2_i), .IN1(na2402_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a433_5 ( .OUT(na433_2), .CLK(na2414_1), .EN(na132_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na433_2_i) );
// C_///AND/D      x139y42     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a434_4 ( .OUT(na434_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a434_5 ( .OUT(na434_2), .CLK(na2414_1), .EN(na132_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na434_2_i) );
// C_AND/D///      x124y48     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a435_1 ( .OUT(na435_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a435_2 ( .OUT(na435_1), .CLK(na2414_1), .EN(na132_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na435_1_i) );
// C_///AND/D      x146y60     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a436_4 ( .OUT(na436_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a436_5 ( .OUT(na436_2), .CLK(na2414_1), .EN(na132_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na436_2_i) );
// C_AND/D///      x150y54     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a437_1 ( .OUT(na437_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a437_2 ( .OUT(na437_1), .CLK(na2414_1), .EN(na132_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na437_1_i) );
// C_AND/D///      x140y62     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a438_1 ( .OUT(na438_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2407_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a438_2 ( .OUT(na438_1), .CLK(na2414_1), .EN(na132_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na438_1_i) );
// C_AND/D///      x139y68     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a439_1 ( .OUT(na439_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a439_2 ( .OUT(na439_1), .CLK(na2414_1), .EN(na132_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na439_1_i) );
// C_///AND/D      x146y80     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a440_4 ( .OUT(na440_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a440_5 ( .OUT(na440_2), .CLK(na2414_1), .EN(na132_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na440_2_i) );
// C_///AND/D      x134y81     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a441_4 ( .OUT(na441_2_i), .IN1(1'b1), .IN2(na2410_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a441_5 ( .OUT(na441_2), .CLK(na2414_1), .EN(na132_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na441_2_i) );
// C_///AND/D      x113y34     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a442_4 ( .OUT(na442_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a442_5 ( .OUT(na442_2), .CLK(na2414_1), .EN(na113_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na442_2_i) );
// C_AND/D///      x106y33     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a443_1 ( .OUT(na443_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a443_2 ( .OUT(na443_1), .CLK(na2414_1), .EN(na113_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na443_1_i) );
// C_AND/D///      x107y44     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a444_1 ( .OUT(na444_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2403_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a444_2 ( .OUT(na444_1), .CLK(na2414_1), .EN(na113_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na444_1_i) );
// C_AND/D///      x105y50     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a445_1 ( .OUT(na445_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a445_2 ( .OUT(na445_1), .CLK(na2414_1), .EN(na113_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na445_1_i) );
// C_///AND/D      x112y58     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a446_4 ( .OUT(na446_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a446_5 ( .OUT(na446_2), .CLK(na2414_1), .EN(na113_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na446_2_i) );
// C_AND/D///      x113y64     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a447_1 ( .OUT(na447_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a447_2 ( .OUT(na447_1), .CLK(na2414_1), .EN(na113_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na447_1_i) );
// C_///AND/D      x109y75     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a448_4 ( .OUT(na448_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a448_5 ( .OUT(na448_2), .CLK(na2414_1), .EN(na113_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na448_2_i) );
// C_///AND/D      x109y79     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a449_4 ( .OUT(na449_2_i), .IN1(na2408_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a449_5 ( .OUT(na449_2), .CLK(na2414_1), .EN(na113_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na449_2_i) );
// C_///AND/D      x114y75     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a450_4 ( .OUT(na450_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a450_5 ( .OUT(na450_2), .CLK(na2414_1), .EN(na113_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na450_2_i) );
// C_AND/D///      x119y78     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a451_1 ( .OUT(na451_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a451_2 ( .OUT(na451_1), .CLK(na2414_1), .EN(na113_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na451_1_i) );
// C_AND/D///      x110y32     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a452_1 ( .OUT(na452_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2401_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a452_2 ( .OUT(na452_1), .CLK(na2414_1), .EN(na99_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na452_1_i) );
// C_AND/D///      x110y38     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a453_1 ( .OUT(na453_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a453_2 ( .OUT(na453_1), .CLK(na2414_1), .EN(na99_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na453_1_i) );
// C_///AND/D      x108y50     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a454_4 ( .OUT(na454_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a454_5 ( .OUT(na454_2), .CLK(na2414_1), .EN(na99_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na454_2_i) );
// C_///AND/D      x111y55     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a455_4 ( .OUT(na455_2_i), .IN1(1'b1), .IN2(na2404_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a455_5 ( .OUT(na455_2), .CLK(na2414_1), .EN(na99_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na455_2_i) );
// C_///AND/D      x112y57     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a456_4 ( .OUT(na456_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a456_5 ( .OUT(na456_2), .CLK(na2414_1), .EN(na99_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na456_2_i) );
// C_AND/D///      x110y60     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a457_1 ( .OUT(na457_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a457_2 ( .OUT(na457_1), .CLK(na2414_1), .EN(na99_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na457_1_i) );
// C_///AND/D      x112y74     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a458_4 ( .OUT(na458_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a458_5 ( .OUT(na458_2), .CLK(na2414_1), .EN(na99_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na458_2_i) );
// C_AND/D///      x110y78     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a459_1 ( .OUT(na459_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a459_2 ( .OUT(na459_1), .CLK(na2414_1), .EN(na99_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na459_1_i) );
// C_AND/D///      x110y79     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a460_1 ( .OUT(na460_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2409_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a460_2 ( .OUT(na460_1), .CLK(na2414_1), .EN(na99_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na460_1_i) );
// C_AND/D///      x120y78     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a461_1 ( .OUT(na461_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a461_2 ( .OUT(na461_1), .CLK(na2414_1), .EN(na99_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na461_1_i) );
// C_///AND/D      x108y33     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a462_4 ( .OUT(na462_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a462_5 ( .OUT(na462_2), .CLK(na2414_1), .EN(na127_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na462_2_i) );
// C_///AND/D      x109y38     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a463_4 ( .OUT(na463_2_i), .IN1(na2402_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a463_5 ( .OUT(na463_2), .CLK(na2414_1), .EN(na127_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na463_2_i) );
// C_///AND/D      x107y48     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a464_4 ( .OUT(na464_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a464_5 ( .OUT(na464_2), .CLK(na2414_1), .EN(na127_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na464_2_i) );
// C_AND/D///      x107y50     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a465_1 ( .OUT(na465_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a465_2 ( .OUT(na465_1), .CLK(na2414_1), .EN(na127_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na465_1_i) );
// C_AND/D///      x105y54     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a466_1 ( .OUT(na466_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2405_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a466_2 ( .OUT(na466_1), .CLK(na2414_1), .EN(na127_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na466_1_i) );
// C_AND/D///      x108y62     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a467_1 ( .OUT(na467_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a467_2 ( .OUT(na467_1), .CLK(na2414_1), .EN(na127_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na467_1_i) );
// C_///AND/D      x107y75     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a468_4 ( .OUT(na468_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a468_5 ( .OUT(na468_2), .CLK(na2414_1), .EN(na127_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na468_2_i) );
// C_AND/D///      x105y80     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a469_1 ( .OUT(na469_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a469_2 ( .OUT(na469_1), .CLK(na2414_1), .EN(na127_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na469_1_i) );
// C_///AND/D      x113y76     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a470_4 ( .OUT(na470_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a470_5 ( .OUT(na470_2), .CLK(na2414_1), .EN(na127_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na470_2_i) );
// C_///AND/D      x127y84     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a471_4 ( .OUT(na471_2_i), .IN1(1'b1), .IN2(na2410_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a471_5 ( .OUT(na471_2), .CLK(na2414_1), .EN(na127_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na471_2_i) );
// C_///AND/D      x109y34     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a472_4 ( .OUT(na472_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a472_5 ( .OUT(na472_2), .CLK(na2414_1), .EN(na126_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na472_2_i) );
// C_AND/D///      x108y37     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a473_1 ( .OUT(na473_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a473_2 ( .OUT(na473_1), .CLK(na2414_1), .EN(na126_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na473_1_i) );
// C_AND/D///      x106y41     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a474_1 ( .OUT(na474_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2403_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a474_2 ( .OUT(na474_1), .CLK(na2414_1), .EN(na126_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na474_1_i) );
// C_AND/D///      x108y49     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a475_1 ( .OUT(na475_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a475_2 ( .OUT(na475_1), .CLK(na2414_1), .EN(na126_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na475_1_i) );
// C_///AND/D      x104y55     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a476_4 ( .OUT(na476_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a476_5 ( .OUT(na476_2), .CLK(na2414_1), .EN(na126_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na476_2_i) );
// C_///AND/D      x109y63     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a477_4 ( .OUT(na477_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2406_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a477_5 ( .OUT(na477_2), .CLK(na2414_1), .EN(na126_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na477_2_i) );
// C_///AND/D      x108y80     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a478_4 ( .OUT(na478_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a478_5 ( .OUT(na478_2), .CLK(na2414_1), .EN(na126_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na478_2_i) );
// C_AND/D///      x108y79     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a479_1 ( .OUT(na479_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a479_2 ( .OUT(na479_1), .CLK(na2414_1), .EN(na126_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na479_1_i) );
// C_///AND/D      x116y73     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a480_4 ( .OUT(na480_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a480_5 ( .OUT(na480_2), .CLK(na2414_1), .EN(na126_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na480_2_i) );
// C_AND/D///      x120y81     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a481_1 ( .OUT(na481_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a481_2 ( .OUT(na481_1), .CLK(na2414_1), .EN(na126_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na481_1_i) );
// C_AND/D///      x105y31     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a482_1 ( .OUT(na482_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2401_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a482_2 ( .OUT(na482_1), .CLK(na2414_1), .EN(na125_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na482_1_i) );
// C_AND/D///      x108y40     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a483_1 ( .OUT(na483_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a483_2 ( .OUT(na483_1), .CLK(na2414_1), .EN(na125_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na483_1_i) );
// C_///AND/D      x112y48     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a484_4 ( .OUT(na484_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a484_5 ( .OUT(na484_2), .CLK(na2414_1), .EN(na125_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na484_2_i) );
// C_///AND/D      x116y56     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a485_4 ( .OUT(na485_2_i), .IN1(1'b1), .IN2(na2404_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a485_5 ( .OUT(na485_2), .CLK(na2414_1), .EN(na125_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na485_2_i) );
// C_///AND/D      x106y54     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a486_4 ( .OUT(na486_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a486_5 ( .OUT(na486_2), .CLK(na2414_1), .EN(na125_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na486_2_i) );
// C_AND/D///      x107y64     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a487_1 ( .OUT(na487_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a487_2 ( .OUT(na487_1), .CLK(na2414_1), .EN(na125_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na487_1_i) );
// C_AND/D///      x108y69     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a488_1 ( .OUT(na488_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2407_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a488_2 ( .OUT(na488_1), .CLK(na2414_1), .EN(na125_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na488_1_i) );
// C_AND/D///      x108y78     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a489_1 ( .OUT(na489_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a489_2 ( .OUT(na489_1), .CLK(na2414_1), .EN(na125_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na489_1_i) );
// C_///AND/D      x114y74     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a490_4 ( .OUT(na490_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a490_5 ( .OUT(na490_2), .CLK(na2414_1), .EN(na125_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na490_2_i) );
// C_AND/D///      x118y82     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a491_1 ( .OUT(na491_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a491_2 ( .OUT(na491_1), .CLK(na2414_1), .EN(na125_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na491_1_i) );
// C_///AND/D      x113y31     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a492_4 ( .OUT(na492_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a492_5 ( .OUT(na492_2), .CLK(na2414_1), .EN(na122_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na492_2_i) );
// C_///AND/D      x109y33     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a493_4 ( .OUT(na493_2_i), .IN1(na2402_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a493_5 ( .OUT(na493_2), .CLK(na2414_1), .EN(na122_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na493_2_i) );
// C_///AND/D      x106y48     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a494_4 ( .OUT(na494_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a494_5 ( .OUT(na494_2), .CLK(na2414_1), .EN(na122_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na494_2_i) );
// C_AND/D///      x108y51     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a495_1 ( .OUT(na495_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a495_2 ( .OUT(na495_1), .CLK(na2414_1), .EN(na122_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na495_1_i) );
// C_AND/D///      x106y55     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a496_1 ( .OUT(na496_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2405_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a496_2 ( .OUT(na496_1), .CLK(na2414_1), .EN(na122_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na496_1_i) );
// C_AND/D///      x108y63     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a497_1 ( .OUT(na497_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a497_2 ( .OUT(na497_1), .CLK(na2414_1), .EN(na122_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na497_1_i) );
// C_///AND/D      x108y73     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a498_4 ( .OUT(na498_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a498_5 ( .OUT(na498_2), .CLK(na2414_1), .EN(na122_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na498_2_i) );
// C_///AND/D      x105y78     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a499_4 ( .OUT(na499_2_i), .IN1(na2408_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a499_5 ( .OUT(na499_2), .CLK(na2414_1), .EN(na122_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na499_2_i) );
// C_///AND/D      x113y80     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a500_4 ( .OUT(na500_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a500_5 ( .OUT(na500_2), .CLK(na2414_1), .EN(na122_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na500_2_i) );
// C_AND/D///      x116y77     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a501_1 ( .OUT(na501_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a501_2 ( .OUT(na501_1), .CLK(na2414_1), .EN(na122_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na501_1_i) );
// C_///AND/D      x106y31     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a502_4 ( .OUT(na502_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a502_5 ( .OUT(na502_2), .CLK(na2414_1), .EN(na103_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na502_2_i) );
// C_AND/D///      x110y37     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a503_1 ( .OUT(na503_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a503_2 ( .OUT(na503_1), .CLK(na2414_1), .EN(na103_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na503_1_i) );
// C_AND/D///      x106y47     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a504_1 ( .OUT(na504_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2403_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a504_2 ( .OUT(na504_1), .CLK(na2414_1), .EN(na103_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na504_1_i) );
// C_AND/D///      x107y54     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a505_1 ( .OUT(na505_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a505_2 ( .OUT(na505_1), .CLK(na2414_1), .EN(na103_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na505_1_i) );
// C_///AND/D      x114y60     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a506_4 ( .OUT(na506_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a506_5 ( .OUT(na506_2), .CLK(na2414_1), .EN(na103_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na506_2_i) );
// C_///AND/D      x110y61     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a507_4 ( .OUT(na507_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2406_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a507_5 ( .OUT(na507_2), .CLK(na2414_1), .EN(na103_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na507_2_i) );
// C_///AND/D      x106y75     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a508_4 ( .OUT(na508_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a508_5 ( .OUT(na508_2), .CLK(na2414_1), .EN(na103_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na508_2_i) );
// C_AND/D///      x106y79     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a509_1 ( .OUT(na509_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a509_2 ( .OUT(na509_1), .CLK(na2414_1), .EN(na103_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na509_1_i) );
// C_AND/D///      x112y84     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a510_1 ( .OUT(na510_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2409_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a510_2 ( .OUT(na510_1), .CLK(na2414_1), .EN(na103_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na510_1_i) );
// C_AND/D///      x120y77     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a511_1 ( .OUT(na511_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a511_2 ( .OUT(na511_1), .CLK(na2414_1), .EN(na103_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na511_1_i) );
// C_///AND/D      x111y34     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a512_4 ( .OUT(na512_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a512_5 ( .OUT(na512_2), .CLK(na2414_1), .EN(na121_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na512_2_i) );
// C_AND/D///      x107y36     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a513_1 ( .OUT(na513_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a513_2 ( .OUT(na513_1), .CLK(na2414_1), .EN(na121_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na513_1_i) );
// C_///AND/D      x106y49     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a514_4 ( .OUT(na514_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a514_5 ( .OUT(na514_2), .CLK(na2414_1), .EN(na121_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na514_2_i) );
// C_///AND/D      x116y54     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a515_4 ( .OUT(na515_2_i), .IN1(1'b1), .IN2(na2404_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a515_5 ( .OUT(na515_2), .CLK(na2414_1), .EN(na121_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na515_2_i) );
// C_///AND/D      x108y52     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a516_4 ( .OUT(na516_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a516_5 ( .OUT(na516_2), .CLK(na2414_1), .EN(na121_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na516_2_i) );
// C_AND/D///      x110y64     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a517_1 ( .OUT(na517_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a517_2 ( .OUT(na517_1), .CLK(na2414_1), .EN(na121_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na517_1_i) );
// C_AND/D///      x110y68     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a518_1 ( .OUT(na518_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2407_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a518_2 ( .OUT(na518_1), .CLK(na2414_1), .EN(na121_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na518_1_i) );
// C_AND/D///      x103y75     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a519_1 ( .OUT(na519_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a519_2 ( .OUT(na519_1), .CLK(na2414_1), .EN(na121_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na519_1_i) );
// C_///AND/D      x113y75     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a520_4 ( .OUT(na520_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a520_5 ( .OUT(na520_2), .CLK(na2414_1), .EN(na121_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na520_2_i) );
// C_///AND/D      x122y82     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a521_4 ( .OUT(na521_2_i), .IN1(1'b1), .IN2(na2410_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a521_5 ( .OUT(na521_2), .CLK(na2414_1), .EN(na121_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na521_2_i) );
// C_///AND/D      x109y32     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a522_4 ( .OUT(na522_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a522_5 ( .OUT(na522_2), .CLK(na2414_1), .EN(na105_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na522_2_i) );
// C_AND/D///      x107y38     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a523_1 ( .OUT(na523_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a523_2 ( .OUT(na523_1), .CLK(na2414_1), .EN(na105_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na523_1_i) );
// C_///AND/D      x109y50     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a524_4 ( .OUT(na524_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a524_5 ( .OUT(na524_2), .CLK(na2414_1), .EN(na105_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na524_2_i) );
// C_AND/D///      x110y53     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a525_1 ( .OUT(na525_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a525_2 ( .OUT(na525_1), .CLK(na2414_1), .EN(na105_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na525_1_i) );
// C_AND/D///      x107y55     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a526_1 ( .OUT(na526_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2405_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a526_2 ( .OUT(na526_1), .CLK(na2414_1), .EN(na105_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na526_1_i) );
// C_AND/D///      x109y62     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a527_1 ( .OUT(na527_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a527_2 ( .OUT(na527_1), .CLK(na2414_1), .EN(na105_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na527_1_i) );
// C_///AND/D      x111y68     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a528_4 ( .OUT(na528_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a528_5 ( .OUT(na528_2), .CLK(na2414_1), .EN(na105_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na528_2_i) );
// C_///AND/D      x107y80     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a529_4 ( .OUT(na529_2_i), .IN1(na2408_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a529_5 ( .OUT(na529_2), .CLK(na2414_1), .EN(na105_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na529_2_i) );
// C_///AND/D      x111y77     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a530_4 ( .OUT(na530_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a530_5 ( .OUT(na530_2), .CLK(na2414_1), .EN(na105_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na530_2_i) );
// C_AND/D///      x117y78     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a531_1 ( .OUT(na531_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a531_2 ( .OUT(na531_1), .CLK(na2414_1), .EN(na105_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na531_1_i) );
// C_AND/D///      x108y31     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a532_1 ( .OUT(na532_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2401_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a532_2 ( .OUT(na532_1), .CLK(na2414_1), .EN(na118_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na532_1_i) );
// C_AND/D///      x110y35     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a533_1 ( .OUT(na533_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a533_2 ( .OUT(na533_1), .CLK(na2414_1), .EN(na118_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na533_1_i) );
// C_///AND/D      x107y52     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a534_4 ( .OUT(na534_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a534_5 ( .OUT(na534_2), .CLK(na2414_1), .EN(na118_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na534_2_i) );
// C_AND/D///      x111y51     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a535_1 ( .OUT(na535_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a535_2 ( .OUT(na535_1), .CLK(na2414_1), .EN(na118_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na535_1_i) );
// C_///AND/D      x109y55     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a536_4 ( .OUT(na536_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a536_5 ( .OUT(na536_2), .CLK(na2414_1), .EN(na118_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na536_2_i) );
// C_///AND/D      x111y61     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a537_4 ( .OUT(na537_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2406_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a537_5 ( .OUT(na537_2), .CLK(na2414_1), .EN(na118_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na537_2_i) );
// C_///AND/D      x109y73     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a538_4 ( .OUT(na538_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a538_5 ( .OUT(na538_2), .CLK(na2414_1), .EN(na118_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na538_2_i) );
// C_AND/D///      x106y78     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a539_1 ( .OUT(na539_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a539_2 ( .OUT(na539_1), .CLK(na2414_1), .EN(na118_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na539_1_i) );
// C_AND/D///      x112y78     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a540_1 ( .OUT(na540_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2409_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a540_2 ( .OUT(na540_1), .CLK(na2414_1), .EN(na118_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na540_1_i) );
// C_AND/D///      x117y77     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a541_1 ( .OUT(na541_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a541_2 ( .OUT(na541_1), .CLK(na2414_1), .EN(na118_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na541_1_i) );
// C_///AND/D      x111y29     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a542_4 ( .OUT(na542_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a542_5 ( .OUT(na542_2), .CLK(na2414_1), .EN(na109_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na542_2_i) );
// C_///AND/D      x109y37     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a543_4 ( .OUT(na543_2_i), .IN1(na2402_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a543_5 ( .OUT(na543_2), .CLK(na2414_1), .EN(na109_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na543_2_i) );
// C_///AND/D      x109y51     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a544_4 ( .OUT(na544_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a544_5 ( .OUT(na544_2), .CLK(na2414_1), .EN(na109_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na544_2_i) );
// C_AND/D///      x110y54     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a545_1 ( .OUT(na545_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a545_2 ( .OUT(na545_1), .CLK(na2414_1), .EN(na109_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na545_1_i) );
// C_///AND/D      x111y60     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a546_4 ( .OUT(na546_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a546_5 ( .OUT(na546_2), .CLK(na2414_1), .EN(na109_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na546_2_i) );
// C_AND/D///      x107y61     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a547_1 ( .OUT(na547_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a547_2 ( .OUT(na547_1), .CLK(na2414_1), .EN(na109_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na547_1_i) );
// C_AND/D///      x111y67     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a548_1 ( .OUT(na548_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2407_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a548_2 ( .OUT(na548_1), .CLK(na2414_1), .EN(na109_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na548_1_i) );
// C_AND/D///      x107y79     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a549_1 ( .OUT(na549_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a549_2 ( .OUT(na549_1), .CLK(na2414_1), .EN(na109_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na549_1_i) );
// C_///AND/D      x111y82     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a550_4 ( .OUT(na550_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a550_5 ( .OUT(na550_2), .CLK(na2414_1), .EN(na109_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na550_2_i) );
// C_///AND/D      x119y79     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a551_4 ( .OUT(na551_2_i), .IN1(1'b1), .IN2(na2410_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a551_5 ( .OUT(na551_2), .CLK(na2414_1), .EN(na109_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na551_2_i) );
// C_///AND/D      x112y34     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a552_4 ( .OUT(na552_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a552_5 ( .OUT(na552_2), .CLK(na2414_1), .EN(na117_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na552_2_i) );
// C_AND/D///      x110y36     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a553_1 ( .OUT(na553_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a553_2 ( .OUT(na553_1), .CLK(na2414_1), .EN(na117_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na553_1_i) );
// C_AND/D///      x105y43     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a554_1 ( .OUT(na554_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2403_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a554_2 ( .OUT(na554_1), .CLK(na2414_1), .EN(na117_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na554_1_i) );
// C_AND/D///      x109y52     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a555_1 ( .OUT(na555_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a555_2 ( .OUT(na555_1), .CLK(na2414_1), .EN(na117_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na555_1_i) );
// C_///AND/D      x107y56     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a556_4 ( .OUT(na556_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a556_5 ( .OUT(na556_2), .CLK(na2414_1), .EN(na117_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na556_2_i) );
// C_AND/D///      x109y64     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a557_1 ( .OUT(na557_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a557_2 ( .OUT(na557_1), .CLK(na2414_1), .EN(na117_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na557_1_i) );
// C_///AND/D      x109y74     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a558_4 ( .OUT(na558_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a558_5 ( .OUT(na558_2), .CLK(na2414_1), .EN(na117_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na558_2_i) );
// C_///AND/D      x104y79     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a559_4 ( .OUT(na559_2_i), .IN1(na2408_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a559_5 ( .OUT(na559_2), .CLK(na2414_1), .EN(na117_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na559_2_i) );
// C_///AND/D      x114y79     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a560_4 ( .OUT(na560_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a560_5 ( .OUT(na560_2), .CLK(na2414_1), .EN(na117_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na560_2_i) );
// C_AND/D///      x117y80     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a561_1 ( .OUT(na561_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a561_2 ( .OUT(na561_1), .CLK(na2414_1), .EN(na117_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na561_1_i) );
// C_AND/D///      x114y32     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a562_1 ( .OUT(na562_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2401_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a562_2 ( .OUT(na562_1), .CLK(na2414_1), .EN(na111_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na562_1_i) );
// C_AND/D///      x107y33     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a563_1 ( .OUT(na563_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a563_2 ( .OUT(na563_1), .CLK(na2414_1), .EN(na111_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na563_1_i) );
// C_///AND/D      x112y50     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a564_4 ( .OUT(na564_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a564_5 ( .OUT(na564_2), .CLK(na2414_1), .EN(na111_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na564_2_i) );
// C_///AND/D      x106y52     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a565_4 ( .OUT(na565_2_i), .IN1(1'b1), .IN2(na2404_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a565_5 ( .OUT(na565_2), .CLK(na2414_1), .EN(na111_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na565_2_i) );
// C_///AND/D      x113y58     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a566_4 ( .OUT(na566_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a566_5 ( .OUT(na566_2), .CLK(na2414_1), .EN(na111_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na566_2_i) );
// C_AND/D///      x114y64     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a567_1 ( .OUT(na567_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a567_2 ( .OUT(na567_1), .CLK(na2414_1), .EN(na111_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na567_1_i) );
// C_///AND/D      x108y77     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a568_4 ( .OUT(na568_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a568_5 ( .OUT(na568_2), .CLK(na2414_1), .EN(na111_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na568_2_i) );
// C_AND/D///      x106y81     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a569_1 ( .OUT(na569_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a569_2 ( .OUT(na569_1), .CLK(na2414_1), .EN(na111_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na569_1_i) );
// C_AND/D///      x113y79     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a570_1 ( .OUT(na570_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2409_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a570_2 ( .OUT(na570_1), .CLK(na2414_1), .EN(na111_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na570_1_i) );
// C_AND/D///      x120y80     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a571_1 ( .OUT(na571_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a571_2 ( .OUT(na571_1), .CLK(na2414_1), .EN(na111_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na571_1_i) );
// C_///AND/D      x113y35     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a572_4 ( .OUT(na572_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a572_5 ( .OUT(na572_2), .CLK(na2414_1), .EN(na114_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na572_2_i) );
// C_///AND/D      x106y36     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a573_4 ( .OUT(na573_2_i), .IN1(na2402_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a573_5 ( .OUT(na573_2), .CLK(na2414_1), .EN(na114_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na573_2_i) );
// C_///AND/D      x113y53     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a574_4 ( .OUT(na574_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a574_5 ( .OUT(na574_2), .CLK(na2414_1), .EN(na114_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na574_2_i) );
// C_AND/D///      x105y51     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a575_1 ( .OUT(na575_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a575_2 ( .OUT(na575_1), .CLK(na2414_1), .EN(na114_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na575_1_i) );
// C_AND/D///      x110y55     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a576_1 ( .OUT(na576_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2405_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a576_2 ( .OUT(na576_1), .CLK(na2414_1), .EN(na114_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na576_1_i) );
// C_AND/D///      x115y63     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a577_1 ( .OUT(na577_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a577_2 ( .OUT(na577_1), .CLK(na2414_1), .EN(na114_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na577_1_i) );
// C_///AND/D      x107y78     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a578_4 ( .OUT(na578_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a578_5 ( .OUT(na578_2), .CLK(na2414_1), .EN(na114_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na578_2_i) );
// C_AND/D///      x107y82     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a579_1 ( .OUT(na579_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a579_2 ( .OUT(na579_1), .CLK(na2414_1), .EN(na114_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na579_1_i) );
// C_///AND/D      x116y80     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a580_4 ( .OUT(na580_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a580_5 ( .OUT(na580_2), .CLK(na2414_1), .EN(na114_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na580_2_i) );
// C_///AND/D      x123y77     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a581_4 ( .OUT(na581_2_i), .IN1(1'b1), .IN2(na2410_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a581_5 ( .OUT(na581_2), .CLK(na2414_1), .EN(na114_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na581_2_i) );
// C_///AND/D      x114y35     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a582_4 ( .OUT(na582_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a582_5 ( .OUT(na582_2), .CLK(na2414_1), .EN(na112_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na582_2_i) );
// C_AND/D///      x105y36     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a583_1 ( .OUT(na583_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a583_2 ( .OUT(na583_1), .CLK(na2414_1), .EN(na112_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na583_1_i) );
// C_AND/D///      x110y45     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a584_1 ( .OUT(na584_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2403_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a584_2 ( .OUT(na584_1), .CLK(na2414_1), .EN(na112_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na584_1_i) );
// C_AND/D///      x110y51     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a585_1 ( .OUT(na585_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a585_2 ( .OUT(na585_1), .CLK(na2414_1), .EN(na112_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na585_1_i) );
// C_///AND/D      x117y57     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a586_4 ( .OUT(na586_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a586_5 ( .OUT(na586_2), .CLK(na2414_1), .EN(na112_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na586_2_i) );
// C_///AND/D      x114y63     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a587_4 ( .OUT(na587_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2406_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a587_5 ( .OUT(na587_2), .CLK(na2414_1), .EN(na112_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na587_2_i) );
// C_///AND/D      x106y80     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a588_4 ( .OUT(na588_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a588_5 ( .OUT(na588_2), .CLK(na2414_1), .EN(na112_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na588_2_i) );
// C_AND/D///      x110y82     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a589_1 ( .OUT(na589_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a589_2 ( .OUT(na589_1), .CLK(na2414_1), .EN(na112_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na589_1_i) );
// C_///AND/D      x117y74     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a590_4 ( .OUT(na590_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a590_5 ( .OUT(na590_2), .CLK(na2414_1), .EN(na112_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na590_2_i) );
// C_AND/D///      x120y79     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a591_1 ( .OUT(na591_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a591_2 ( .OUT(na591_1), .CLK(na2414_1), .EN(na112_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na591_1_i) );
// C_AND/D///      x150y38     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a592_1 ( .OUT(na592_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2401_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a592_2 ( .OUT(na592_1), .CLK(na2414_1), .EN(na81_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na592_1_i) );
// C_AND/D///      x139y32     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a593_1 ( .OUT(na593_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a593_2 ( .OUT(na593_1), .CLK(na2414_1), .EN(na81_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na593_1_i) );
// C_///AND/D      x135y43     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a594_4 ( .OUT(na594_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a594_5 ( .OUT(na594_2), .CLK(na2414_1), .EN(na81_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na594_2_i) );
// C_///AND/D      x126y48     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a595_4 ( .OUT(na595_2_i), .IN1(1'b1), .IN2(na2404_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a595_5 ( .OUT(na595_2), .CLK(na2414_1), .EN(na81_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na595_2_i) );
// C_///AND/D      x147y59     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a596_4 ( .OUT(na596_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a596_5 ( .OUT(na596_2), .CLK(na2414_1), .EN(na81_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na596_2_i) );
// C_AND/D///      x146y50     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a597_1 ( .OUT(na597_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a597_2 ( .OUT(na597_1), .CLK(na2414_1), .EN(na81_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na597_1_i) );
// C_AND/D///      x144y64     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a598_1 ( .OUT(na598_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2407_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a598_2 ( .OUT(na598_1), .CLK(na2414_1), .EN(na81_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na598_1_i) );
// C_AND/D///      x140y66     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a599_1 ( .OUT(na599_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a599_2 ( .OUT(na599_1), .CLK(na2414_1), .EN(na81_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na599_1_i) );
// C_///AND/D      x139y75     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a600_4 ( .OUT(na600_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a600_5 ( .OUT(na600_2), .CLK(na2414_1), .EN(na81_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na600_2_i) );
// C_AND/D///      x125y82     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a601_1 ( .OUT(na601_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a601_2 ( .OUT(na601_1), .CLK(na2414_1), .EN(na81_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na601_1_i) );
// C_///AND/D      x146y34     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a602_4 ( .OUT(na602_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a602_5 ( .OUT(na602_2), .CLK(na2414_1), .EN(na150_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na602_2_i) );
// C_///AND/D      x147y35     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a603_4 ( .OUT(na603_2_i), .IN1(na2402_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a603_5 ( .OUT(na603_2), .CLK(na2414_1), .EN(na150_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na603_2_i) );
// C_///AND/D      x141y58     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a604_4 ( .OUT(na604_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a604_5 ( .OUT(na604_2), .CLK(na2414_1), .EN(na150_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na604_2_i) );
// C_AND/D///      x132y54     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a605_1 ( .OUT(na605_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a605_2 ( .OUT(na605_1), .CLK(na2414_1), .EN(na150_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na605_1_i) );
// C_AND/D///      x154y41     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a606_1 ( .OUT(na606_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2405_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a606_2 ( .OUT(na606_1), .CLK(na2414_1), .EN(na150_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na606_1_i) );
// C_AND/D///      x150y53     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a607_1 ( .OUT(na607_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a607_2 ( .OUT(na607_1), .CLK(na2414_1), .EN(na150_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na607_1_i) );
// C_///AND/D      x144y60     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a608_4 ( .OUT(na608_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a608_5 ( .OUT(na608_2), .CLK(na2414_1), .EN(na150_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na608_2_i) );
// C_///AND/D      x140y74     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a609_4 ( .OUT(na609_2_i), .IN1(na2408_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a609_5 ( .OUT(na609_2), .CLK(na2414_1), .EN(na150_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na609_2_i) );
// C_///AND/D      x150y81     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a610_4 ( .OUT(na610_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a610_5 ( .OUT(na610_2), .CLK(na2414_1), .EN(na150_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na610_2_i) );
// C_AND/D///      x136y84     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a611_1 ( .OUT(na611_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a611_2 ( .OUT(na611_1), .CLK(na2414_1), .EN(na150_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na611_1_i) );
// C_///AND/D      x143y34     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a612_4 ( .OUT(na612_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a612_5 ( .OUT(na612_2), .CLK(na2414_1), .EN(na136_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na612_2_i) );
// C_AND/D///      x146y32     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a613_1 ( .OUT(na613_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a613_2 ( .OUT(na613_1), .CLK(na2414_1), .EN(na136_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na613_1_i) );
// C_AND/D///      x145y42     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a614_1 ( .OUT(na614_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2403_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a614_2 ( .OUT(na614_1), .CLK(na2414_1), .EN(na136_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na614_1_i) );
// C_AND/D///      x129y50     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a615_1 ( .OUT(na615_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a615_2 ( .OUT(na615_1), .CLK(na2414_1), .EN(na136_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na615_1_i) );
// C_///AND/D      x151y47     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a616_4 ( .OUT(na616_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a616_5 ( .OUT(na616_2), .CLK(na2414_1), .EN(na136_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na616_2_i) );
// C_///AND/D      x147y62     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a617_4 ( .OUT(na617_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2406_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a617_5 ( .OUT(na617_2), .CLK(na2414_1), .EN(na136_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na617_2_i) );
// C_///AND/D      x135y62     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a618_4 ( .OUT(na618_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a618_5 ( .OUT(na618_2), .CLK(na2414_1), .EN(na136_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na618_2_i) );
// C_AND/D///      x145y73     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a619_1 ( .OUT(na619_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a619_2 ( .OUT(na619_1), .CLK(na2414_1), .EN(na136_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na619_1_i) );
// C_AND/D///      x150y78     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a620_1 ( .OUT(na620_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2409_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a620_2 ( .OUT(na620_1), .CLK(na2414_1), .EN(na136_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na620_1_i) );
// C_AND/D///      x135y79     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a621_1 ( .OUT(na621_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a621_2 ( .OUT(na621_1), .CLK(na2414_1), .EN(na136_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na621_1_i) );
// C_///AND/D      x144y35     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a622_4 ( .OUT(na622_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a622_5 ( .OUT(na622_2), .CLK(na2414_1), .EN(na137_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na622_2_i) );
// C_AND/D///      x143y31     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a623_1 ( .OUT(na623_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a623_2 ( .OUT(na623_1), .CLK(na2414_1), .EN(na137_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na623_1_i) );
// C_///AND/D      x144y49     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a624_4 ( .OUT(na624_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a624_5 ( .OUT(na624_2), .CLK(na2414_1), .EN(na137_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na624_2_i) );
// C_///AND/D      x134y45     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a625_4 ( .OUT(na625_2_i), .IN1(1'b1), .IN2(na2404_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a625_5 ( .OUT(na625_2), .CLK(na2414_1), .EN(na137_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na625_2_i) );
// C_///AND/D      x156y46     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a626_4 ( .OUT(na626_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a626_5 ( .OUT(na626_2), .CLK(na2414_1), .EN(na137_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na626_2_i) );
// C_AND/D///      x150y49     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a627_1 ( .OUT(na627_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a627_2 ( .OUT(na627_1), .CLK(na2414_1), .EN(na137_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na627_1_i) );
// C_AND/D///      x146y63     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a628_1 ( .OUT(na628_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2407_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a628_2 ( .OUT(na628_1), .CLK(na2414_1), .EN(na137_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na628_1_i) );
// C_AND/D///      x150y74     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a629_1 ( .OUT(na629_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a629_2 ( .OUT(na629_1), .CLK(na2414_1), .EN(na137_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na629_1_i) );
// C_///AND/D      x149y75     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a630_4 ( .OUT(na630_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a630_5 ( .OUT(na630_2), .CLK(na2414_1), .EN(na137_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na630_2_i) );
// C_///AND/D      x138y84     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a631_4 ( .OUT(na631_2_i), .IN1(1'b1), .IN2(na2410_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a631_5 ( .OUT(na631_2), .CLK(na2414_1), .EN(na137_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na631_2_i) );
// C_///AND/D      x144y34     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a632_4 ( .OUT(na632_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a632_5 ( .OUT(na632_2), .CLK(na2414_1), .EN(na138_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na632_2_i) );
// C_AND/D///      x145y32     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a633_1 ( .OUT(na633_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a633_2 ( .OUT(na633_1), .CLK(na2414_1), .EN(na138_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na633_1_i) );
// C_///AND/D      x142y52     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a634_4 ( .OUT(na634_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a634_5 ( .OUT(na634_2), .CLK(na2414_1), .EN(na138_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na634_2_i) );
// C_AND/D///      x128y50     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a635_1 ( .OUT(na635_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a635_2 ( .OUT(na635_1), .CLK(na2414_1), .EN(na138_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na635_1_i) );
// C_AND/D///      x154y39     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a636_1 ( .OUT(na636_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2405_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a636_2 ( .OUT(na636_1), .CLK(na2414_1), .EN(na138_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na636_1_i) );
// C_AND/D///      x152y52     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a637_1 ( .OUT(na637_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a637_2 ( .OUT(na637_1), .CLK(na2414_1), .EN(na138_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na637_1_i) );
// C_///AND/D      x136y64     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a638_4 ( .OUT(na638_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a638_5 ( .OUT(na638_2), .CLK(na2414_1), .EN(na138_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na638_2_i) );
// C_///AND/D      x144y77     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a639_4 ( .OUT(na639_2_i), .IN1(na2408_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a639_5 ( .OUT(na639_2), .CLK(na2414_1), .EN(na138_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na639_2_i) );
// C_///AND/D      x151y74     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a640_4 ( .OUT(na640_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a640_5 ( .OUT(na640_2), .CLK(na2414_1), .EN(na138_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na640_2_i) );
// C_AND/D///      x136y79     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a641_1 ( .OUT(na641_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a641_2 ( .OUT(na641_1), .CLK(na2414_1), .EN(na138_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na641_1_i) );
// C_AND/D///      x145y35     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a642_1 ( .OUT(na642_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2401_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a642_2 ( .OUT(na642_1), .CLK(na2414_1), .EN(na139_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na642_1_i) );
// C_AND/D///      x148y31     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a643_1 ( .OUT(na643_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a643_2 ( .OUT(na643_1), .CLK(na2414_1), .EN(na139_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na643_1_i) );
// C_///AND/D      x144y50     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a644_4 ( .OUT(na644_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a644_5 ( .OUT(na644_2), .CLK(na2414_1), .EN(na139_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na644_2_i) );
// C_AND/D///      x129y52     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a645_1 ( .OUT(na645_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a645_2 ( .OUT(na645_1), .CLK(na2414_1), .EN(na139_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na645_1_i) );
// C_///AND/D      x153y52     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a646_4 ( .OUT(na646_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a646_5 ( .OUT(na646_2), .CLK(na2414_1), .EN(na139_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na646_2_i) );
// C_///AND/D      x145y57     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a647_4 ( .OUT(na647_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2406_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a647_5 ( .OUT(na647_2), .CLK(na2414_1), .EN(na139_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na647_2_i) );
// C_///AND/D      x141y68     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a648_4 ( .OUT(na648_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a648_5 ( .OUT(na648_2), .CLK(na2414_1), .EN(na139_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na648_2_i) );
// C_AND/D///      x148y70     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a649_1 ( .OUT(na649_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a649_2 ( .OUT(na649_1), .CLK(na2414_1), .EN(na139_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na649_1_i) );
// C_AND/D///      x152y74     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a650_1 ( .OUT(na650_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2409_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a650_2 ( .OUT(na650_1), .CLK(na2414_1), .EN(na139_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na650_1_i) );
// C_AND/D///      x131y83     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a651_1 ( .OUT(na651_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a651_2 ( .OUT(na651_1), .CLK(na2414_1), .EN(na139_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na651_1_i) );
// C_///AND/D      x145y36     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a652_4 ( .OUT(na652_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a652_5 ( .OUT(na652_2), .CLK(na2414_1), .EN(na140_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na652_2_i) );
// C_///AND/D      x148y34     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a653_4 ( .OUT(na653_2_i), .IN1(na2402_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a653_5 ( .OUT(na653_2), .CLK(na2414_1), .EN(na140_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na653_2_i) );
// C_///AND/D      x148y49     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a654_4 ( .OUT(na654_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a654_5 ( .OUT(na654_2), .CLK(na2414_1), .EN(na140_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na654_2_i) );
// C_AND/D///      x127y51     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a655_1 ( .OUT(na655_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a655_2 ( .OUT(na655_1), .CLK(na2414_1), .EN(na140_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na655_1_i) );
// C_///AND/D      x153y49     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a656_4 ( .OUT(na656_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a656_5 ( .OUT(na656_2), .CLK(na2414_1), .EN(na140_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na656_2_i) );
// C_AND/D///      x145y52     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a657_1 ( .OUT(na657_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a657_2 ( .OUT(na657_1), .CLK(na2414_1), .EN(na140_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na657_1_i) );
// C_AND/D///      x143y61     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a658_1 ( .OUT(na658_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2407_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a658_2 ( .OUT(na658_1), .CLK(na2414_1), .EN(na140_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na658_1_i) );
// C_AND/D///      x146y71     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a659_1 ( .OUT(na659_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a659_2 ( .OUT(na659_1), .CLK(na2414_1), .EN(na140_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na659_1_i) );
// C_///AND/D      x152y77     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a660_4 ( .OUT(na660_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a660_5 ( .OUT(na660_2), .CLK(na2414_1), .EN(na140_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na660_2_i) );
// C_///AND/D      x137y84     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a661_4 ( .OUT(na661_2_i), .IN1(1'b1), .IN2(na2410_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a661_5 ( .OUT(na661_2), .CLK(na2414_1), .EN(na140_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na661_2_i) );
// C_///AND/D      x144y37     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a662_4 ( .OUT(na662_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a662_5 ( .OUT(na662_2), .CLK(na2414_1), .EN(na141_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na662_2_i) );
// C_AND/D///      x149y33     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a663_1 ( .OUT(na663_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a663_2 ( .OUT(na663_1), .CLK(na2414_1), .EN(na141_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na663_1_i) );
// C_AND/D///      x149y42     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a664_1 ( .OUT(na664_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2403_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a664_2 ( .OUT(na664_1), .CLK(na2414_1), .EN(na141_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na664_1_i) );
// C_AND/D///      x130y52     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a665_1 ( .OUT(na665_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a665_2 ( .OUT(na665_1), .CLK(na2414_1), .EN(na141_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na665_1_i) );
// C_///AND/D      x156y52     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a666_4 ( .OUT(na666_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a666_5 ( .OUT(na666_2), .CLK(na2414_1), .EN(na141_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na666_2_i) );
// C_AND/D///      x150y51     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a667_1 ( .OUT(na667_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a667_2 ( .OUT(na667_1), .CLK(na2414_1), .EN(na141_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na667_1_i) );
// C_///AND/D      x142y68     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a668_4 ( .OUT(na668_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a668_5 ( .OUT(na668_2), .CLK(na2414_1), .EN(na141_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na668_2_i) );
// C_///AND/D      x143y76     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a669_4 ( .OUT(na669_2_i), .IN1(na2408_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a669_5 ( .OUT(na669_2), .CLK(na2414_1), .EN(na141_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na669_2_i) );
// C_///AND/D      x147y80     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a670_4 ( .OUT(na670_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a670_5 ( .OUT(na670_2), .CLK(na2414_1), .EN(na141_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na670_2_i) );
// C_AND/D///      x132y81     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a671_1 ( .OUT(na671_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a671_2 ( .OUT(na671_1), .CLK(na2414_1), .EN(na141_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na671_1_i) );
// C_AND/D///      x150y34     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a672_1 ( .OUT(na672_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2401_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a672_2 ( .OUT(na672_1), .CLK(na2414_1), .EN(na142_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na672_1_i) );
// C_AND/D///      x149y32     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a673_1 ( .OUT(na673_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a673_2 ( .OUT(na673_1), .CLK(na2414_1), .EN(na142_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na673_1_i) );
// C_///AND/D      x147y51     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a674_4 ( .OUT(na674_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a674_5 ( .OUT(na674_2), .CLK(na2414_1), .EN(na142_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na674_2_i) );
// C_///AND/D      x126y49     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a675_4 ( .OUT(na675_2_i), .IN1(1'b1), .IN2(na2404_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a675_5 ( .OUT(na675_2), .CLK(na2414_1), .EN(na142_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na675_2_i) );
// C_///AND/D      x156y51     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a676_4 ( .OUT(na676_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a676_5 ( .OUT(na676_2), .CLK(na2414_1), .EN(na142_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na676_2_i) );
// C_AND/D///      x148y52     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a677_1 ( .OUT(na677_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a677_2 ( .OUT(na677_1), .CLK(na2414_1), .EN(na142_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na677_1_i) );
// C_///AND/D      x142y69     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a678_4 ( .OUT(na678_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a678_5 ( .OUT(na678_2), .CLK(na2414_1), .EN(na142_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na678_2_i) );
// C_AND/D///      x147y71     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a679_1 ( .OUT(na679_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a679_2 ( .OUT(na679_1), .CLK(na2414_1), .EN(na142_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na679_1_i) );
// C_AND/D///      x151y75     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a680_1 ( .OUT(na680_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2409_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a680_2 ( .OUT(na680_1), .CLK(na2414_1), .EN(na142_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na680_1_i) );
// C_AND/D///      x134y82     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a681_1 ( .OUT(na681_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a681_2 ( .OUT(na681_1), .CLK(na2414_1), .EN(na142_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na681_1_i) );
// C_///AND/D      x143y37     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a682_4 ( .OUT(na682_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a682_5 ( .OUT(na682_2), .CLK(na2414_1), .EN(na143_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na682_2_i) );
// C_///AND/D      x147y33     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a683_4 ( .OUT(na683_2_i), .IN1(na2402_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a683_5 ( .OUT(na683_2), .CLK(na2414_1), .EN(na143_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na683_2_i) );
// C_///AND/D      x142y42     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a684_4 ( .OUT(na684_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a684_5 ( .OUT(na684_2), .CLK(na2414_1), .EN(na143_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na684_2_i) );
// C_AND/D///      x131y50     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a685_1 ( .OUT(na685_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a685_2 ( .OUT(na685_1), .CLK(na2414_1), .EN(na143_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na685_1_i) );
// C_AND/D///      x154y43     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a686_1 ( .OUT(na686_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2405_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a686_2 ( .OUT(na686_1), .CLK(na2414_1), .EN(na143_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na686_1_i) );
// C_AND/D///      x155y49     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a687_1 ( .OUT(na687_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a687_2 ( .OUT(na687_1), .CLK(na2414_1), .EN(na143_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na687_1_i) );
// C_///AND/D      x141y61     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a688_4 ( .OUT(na688_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a688_5 ( .OUT(na688_2), .CLK(na2414_1), .EN(na143_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na688_2_i) );
// C_AND/D///      x143y70     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a689_1 ( .OUT(na689_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a689_2 ( .OUT(na689_1), .CLK(na2414_1), .EN(na143_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na689_1_i) );
// C_///AND/D      x148y79     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a690_4 ( .OUT(na690_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a690_5 ( .OUT(na690_2), .CLK(na2414_1), .EN(na143_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na690_2_i) );
// C_///AND/D      x139y81     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a691_4 ( .OUT(na691_2_i), .IN1(1'b1), .IN2(na2410_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a691_5 ( .OUT(na691_2), .CLK(na2414_1), .EN(na143_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na691_2_i) );
// C_///AND/D      x143y35     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a692_4 ( .OUT(na692_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a692_5 ( .OUT(na692_2), .CLK(na2414_1), .EN(na133_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na692_2_i) );
// C_AND/D///      x146y29     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a693_1 ( .OUT(na693_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a693_2 ( .OUT(na693_1), .CLK(na2414_1), .EN(na133_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na693_1_i) );
// C_AND/D///      x147y41     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a694_1 ( .OUT(na694_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2403_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a694_2 ( .OUT(na694_1), .CLK(na2414_1), .EN(na133_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na694_1_i) );
// C_AND/D///      x129y49     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a695_1 ( .OUT(na695_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a695_2 ( .OUT(na695_1), .CLK(na2414_1), .EN(na133_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na695_1_i) );
// C_///AND/D      x155y48     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a696_4 ( .OUT(na696_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a696_5 ( .OUT(na696_2), .CLK(na2414_1), .EN(na133_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na696_2_i) );
// C_///AND/D      x147y63     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a697_4 ( .OUT(na697_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2406_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a697_5 ( .OUT(na697_2), .CLK(na2414_1), .EN(na133_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na697_2_i) );
// C_///AND/D      x139y63     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a698_4 ( .OUT(na698_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a698_5 ( .OUT(na698_2), .CLK(na2414_1), .EN(na133_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na698_2_i) );
// C_AND/D///      x147y76     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a699_1 ( .OUT(na699_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a699_2 ( .OUT(na699_1), .CLK(na2414_1), .EN(na133_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na699_1_i) );
// C_///AND/D      x156y67     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a700_4 ( .OUT(na700_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a700_5 ( .OUT(na700_2), .CLK(na2414_1), .EN(na133_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na700_2_i) );
// C_AND/D///      x135y80     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a701_1 ( .OUT(na701_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a701_2 ( .OUT(na701_1), .CLK(na2414_1), .EN(na133_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na701_1_i) );
// C_AND/D///      x150y35     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a702_1 ( .OUT(na702_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2401_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a702_2 ( .OUT(na702_1), .CLK(na2414_1), .EN(na145_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na702_1_i) );
// C_AND/D///      x154y31     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a703_1 ( .OUT(na703_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a703_2 ( .OUT(na703_1), .CLK(na2414_1), .EN(na145_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na703_1_i) );
// C_///AND/D      x137y44     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a704_4 ( .OUT(na704_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a704_5 ( .OUT(na704_2), .CLK(na2414_1), .EN(na145_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na704_2_i) );
// C_///AND/D      x136y46     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a705_4 ( .OUT(na705_2_i), .IN1(1'b1), .IN2(na2404_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a705_5 ( .OUT(na705_2), .CLK(na2414_1), .EN(na145_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na705_2_i) );
// C_///AND/D      x149y51     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a706_4 ( .OUT(na706_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a706_5 ( .OUT(na706_2), .CLK(na2414_1), .EN(na145_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na706_2_i) );
// C_AND/D///      x154y51     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a707_1 ( .OUT(na707_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a707_2 ( .OUT(na707_1), .CLK(na2414_1), .EN(na145_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na707_1_i) );
// C_AND/D///      x148y63     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a708_1 ( .OUT(na708_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2407_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a708_2 ( .OUT(na708_1), .CLK(na2414_1), .EN(na145_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na708_1_i) );
// C_AND/D///      x144y72     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a709_1 ( .OUT(na709_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a709_2 ( .OUT(na709_1), .CLK(na2414_1), .EN(na145_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na709_1_i) );
// C_///AND/D      x149y79     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a710_4 ( .OUT(na710_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a710_5 ( .OUT(na710_2), .CLK(na2414_1), .EN(na145_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na710_2_i) );
// C_AND/D///      x138y77     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a711_1 ( .OUT(na711_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a711_2 ( .OUT(na711_1), .CLK(na2414_1), .EN(na145_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na711_1_i) );
// C_///AND/D      x142y38     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a712_4 ( .OUT(na712_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a712_5 ( .OUT(na712_2), .CLK(na2414_1), .EN(na146_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na712_2_i) );
// C_///AND/D      x154y34     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a713_4 ( .OUT(na713_2_i), .IN1(na2402_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a713_5 ( .OUT(na713_2), .CLK(na2414_1), .EN(na146_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na713_2_i) );
// C_///AND/D      x141y47     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a714_4 ( .OUT(na714_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a714_5 ( .OUT(na714_2), .CLK(na2414_1), .EN(na146_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na714_2_i) );
// C_AND/D///      x134y49     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a715_1 ( .OUT(na715_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a715_2 ( .OUT(na715_1), .CLK(na2414_1), .EN(na146_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na715_1_i) );
// C_AND/D///      x153y44     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a716_1 ( .OUT(na716_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2405_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a716_2 ( .OUT(na716_1), .CLK(na2414_1), .EN(na146_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na716_1_i) );
// C_AND/D///      x154y52     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a717_1 ( .OUT(na717_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a717_2 ( .OUT(na717_1), .CLK(na2414_1), .EN(na146_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na717_1_i) );
// C_///AND/D      x142y64     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a718_4 ( .OUT(na718_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a718_5 ( .OUT(na718_2), .CLK(na2414_1), .EN(na146_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na718_2_i) );
// C_///AND/D      x142y77     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a719_4 ( .OUT(na719_2_i), .IN1(na2408_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a719_5 ( .OUT(na719_2), .CLK(na2414_1), .EN(na146_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na719_2_i) );
// C_///AND/D      x143y82     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a720_4 ( .OUT(na720_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a720_5 ( .OUT(na720_2), .CLK(na2414_1), .EN(na146_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na720_2_i) );
// C_AND/D///      x134y80     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a721_1 ( .OUT(na721_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a721_2 ( .OUT(na721_1), .CLK(na2414_1), .EN(na146_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na721_1_i) );
// C_///AND/D      x141y35     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a722_4 ( .OUT(na722_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a722_5 ( .OUT(na722_2), .CLK(na2414_1), .EN(na147_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na722_2_i) );
// C_AND/D///      x150y32     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a723_1 ( .OUT(na723_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a723_2 ( .OUT(na723_1), .CLK(na2414_1), .EN(na147_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na723_1_i) );
// C_AND/D///      x148y43     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a724_1 ( .OUT(na724_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2403_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a724_2 ( .OUT(na724_1), .CLK(na2414_1), .EN(na147_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na724_1_i) );
// C_AND/D///      x131y55     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a725_1 ( .OUT(na725_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a725_2 ( .OUT(na725_1), .CLK(na2414_1), .EN(na147_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na725_1_i) );
// C_///AND/D      x145y54     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a726_4 ( .OUT(na726_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a726_5 ( .OUT(na726_2), .CLK(na2414_1), .EN(na147_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na726_2_i) );
// C_///AND/D      x145y62     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a727_4 ( .OUT(na727_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2406_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a727_5 ( .OUT(na727_2), .CLK(na2414_1), .EN(na147_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na727_2_i) );
// C_///AND/D      x141y63     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a728_4 ( .OUT(na728_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a728_5 ( .OUT(na728_2), .CLK(na2414_1), .EN(na147_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na728_2_i) );
// C_AND/D///      x145y71     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a729_1 ( .OUT(na729_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a729_2 ( .OUT(na729_1), .CLK(na2414_1), .EN(na147_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na729_1_i) );
// C_AND/D///      x151y80     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a730_1 ( .OUT(na730_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2409_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a730_2 ( .OUT(na730_1), .CLK(na2414_1), .EN(na147_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na730_1_i) );
// C_AND/D///      x137y81     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a731_1 ( .OUT(na731_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a731_2 ( .OUT(na731_1), .CLK(na2414_1), .EN(na147_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na731_1_i) );
// C_///AND/D      x143y40     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a732_4 ( .OUT(na732_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a732_5 ( .OUT(na732_2), .CLK(na2414_1), .EN(na148_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na732_2_i) );
// C_AND/D///      x152y31     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a733_1 ( .OUT(na733_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a733_2 ( .OUT(na733_1), .CLK(na2414_1), .EN(na148_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na733_1_i) );
// C_///AND/D      x146y54     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a734_4 ( .OUT(na734_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a734_5 ( .OUT(na734_2), .CLK(na2414_1), .EN(na148_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na734_2_i) );
// C_///AND/D      x127y50     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a735_4 ( .OUT(na735_2_i), .IN1(1'b1), .IN2(na2404_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a735_5 ( .OUT(na735_2), .CLK(na2414_1), .EN(na148_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na735_2_i) );
// C_///AND/D      x149y53     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a736_4 ( .OUT(na736_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a736_5 ( .OUT(na736_2), .CLK(na2414_1), .EN(na148_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na736_2_i) );
// C_AND/D///      x149y53     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a737_1 ( .OUT(na737_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a737_2 ( .OUT(na737_1), .CLK(na2414_1), .EN(na148_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na737_1_i) );
// C_AND/D///      x149y62     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a738_1 ( .OUT(na738_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2407_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a738_2 ( .OUT(na738_1), .CLK(na2414_1), .EN(na148_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na738_1_i) );
// C_AND/D///      x145y76     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a739_1 ( .OUT(na739_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a739_2 ( .OUT(na739_1), .CLK(na2414_1), .EN(na148_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na739_1_i) );
// C_///AND/D      x149y71     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a740_4 ( .OUT(na740_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a740_5 ( .OUT(na740_2), .CLK(na2414_1), .EN(na148_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na740_2_i) );
// C_///AND/D      x139y84     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a741_4 ( .OUT(na741_2_i), .IN1(1'b1), .IN2(na2410_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a741_5 ( .OUT(na741_2), .CLK(na2414_1), .EN(na148_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na741_2_i) );
// C_///AND/D      x146y39     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a742_4 ( .OUT(na742_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a742_5 ( .OUT(na742_2), .CLK(na2414_1), .EN(na149_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na742_2_i) );
// C_AND/D///      x151y32     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a743_1 ( .OUT(na743_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a743_2 ( .OUT(na743_1), .CLK(na2414_1), .EN(na149_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na743_1_i) );
// C_///AND/D      x143y55     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a744_4 ( .OUT(na744_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a744_5 ( .OUT(na744_2), .CLK(na2414_1), .EN(na149_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na744_2_i) );
// C_AND/D///      x132y55     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a745_1 ( .OUT(na745_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a745_2 ( .OUT(na745_1), .CLK(na2414_1), .EN(na149_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na745_1_i) );
// C_AND/D///      x152y42     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a746_1 ( .OUT(na746_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2405_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a746_2 ( .OUT(na746_1), .CLK(na2414_1), .EN(na149_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na746_1_i) );
// C_AND/D///      x152y54     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a747_1 ( .OUT(na747_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a747_2 ( .OUT(na747_1), .CLK(na2414_1), .EN(na149_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na747_1_i) );
// C_///AND/D      x142y61     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a748_4 ( .OUT(na748_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a748_5 ( .OUT(na748_2), .CLK(na2414_1), .EN(na149_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na748_2_i) );
// C_///AND/D      x146y75     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a749_4 ( .OUT(na749_2_i), .IN1(na2408_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a749_5 ( .OUT(na749_2), .CLK(na2414_1), .EN(na149_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na749_2_i) );
// C_///AND/D      x152y78     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a750_4 ( .OUT(na750_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a750_5 ( .OUT(na750_2), .CLK(na2414_1), .EN(na149_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na750_2_i) );
// C_AND/D///      x138y81     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a751_1 ( .OUT(na751_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a751_2 ( .OUT(na751_1), .CLK(na2414_1), .EN(na149_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na751_1_i) );
// C_AND/D///      x149y36     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a752_1 ( .OUT(na752_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2401_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a752_2 ( .OUT(na752_1), .CLK(na2414_1), .EN(na144_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na752_1_i) );
// C_AND/D///      x153y32     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a753_1 ( .OUT(na753_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a753_2 ( .OUT(na753_1), .CLK(na2414_1), .EN(na144_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na753_1_i) );
// C_///AND/D      x134y43     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a754_4 ( .OUT(na754_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a754_5 ( .OUT(na754_2), .CLK(na2414_1), .EN(na144_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na754_2_i) );
// C_AND/D///      x133y51     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a755_1 ( .OUT(na755_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a755_2 ( .OUT(na755_1), .CLK(na2414_1), .EN(na144_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na755_1_i) );
// C_///AND/D      x156y54     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a756_4 ( .OUT(na756_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a756_5 ( .OUT(na756_2), .CLK(na2414_1), .EN(na144_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na756_2_i) );
// C_///AND/D      x153y64     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a757_4 ( .OUT(na757_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2406_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a757_5 ( .OUT(na757_2), .CLK(na2414_1), .EN(na144_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na757_2_i) );
// C_///AND/D      x143y66     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a758_4 ( .OUT(na758_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a758_5 ( .OUT(na758_2), .CLK(na2414_1), .EN(na144_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na758_2_i) );
// C_AND/D///      x143y71     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a759_1 ( .OUT(na759_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a759_2 ( .OUT(na759_1), .CLK(na2414_1), .EN(na144_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na759_1_i) );
// C_AND/D///      x150y80     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a760_1 ( .OUT(na760_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2409_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a760_2 ( .OUT(na760_1), .CLK(na2414_1), .EN(na144_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na760_1_i) );
// C_AND/D///      x137y80     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a761_1 ( .OUT(na761_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a761_2 ( .OUT(na761_1), .CLK(na2414_1), .EN(na144_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na761_1_i) );
// C_///AND/D      x121y31     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a762_4 ( .OUT(na762_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a762_5 ( .OUT(na762_2), .CLK(na2414_1), .EN(na168_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na762_2_i) );
// C_///AND/D      x124y42     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a763_4 ( .OUT(na763_2_i), .IN1(na2402_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a763_5 ( .OUT(na763_2), .CLK(na2414_1), .EN(na168_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na763_2_i) );
// C_///AND/D      x116y41     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a764_4 ( .OUT(na764_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a764_5 ( .OUT(na764_2), .CLK(na2414_1), .EN(na168_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na764_2_i) );
// C_AND/D///      x120y44     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a765_1 ( .OUT(na765_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a765_2 ( .OUT(na765_1), .CLK(na2414_1), .EN(na168_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na765_1_i) );
// C_///AND/D      x118y53     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a766_4 ( .OUT(na766_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a766_5 ( .OUT(na766_2), .CLK(na2414_1), .EN(na168_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na766_2_i) );
// C_AND/D///      x128y53     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a767_1 ( .OUT(na767_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a767_2 ( .OUT(na767_1), .CLK(na2414_1), .EN(na168_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na767_1_i) );
// C_AND/D///      x129y66     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a768_1 ( .OUT(na768_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2407_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a768_2 ( .OUT(na768_1), .CLK(na2414_1), .EN(na168_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na768_1_i) );
// C_AND/D///      x122y69     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a769_1 ( .OUT(na769_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a769_2 ( .OUT(na769_1), .CLK(na2414_1), .EN(na168_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na769_1_i) );
// C_///AND/D      x118y78     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a770_4 ( .OUT(na770_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a770_5 ( .OUT(na770_2), .CLK(na2414_1), .EN(na168_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na770_2_i) );
// C_///AND/D      x129y79     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a771_4 ( .OUT(na771_2_i), .IN1(1'b1), .IN2(na2410_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a771_5 ( .OUT(na771_2), .CLK(na2414_1), .EN(na168_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na771_2_i) );
// C_///AND/D      x115y31     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a772_4 ( .OUT(na772_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a772_5 ( .OUT(na772_2), .CLK(na2414_1), .EN(na154_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na772_2_i) );
// C_AND/D///      x117y34     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a773_1 ( .OUT(na773_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a773_2 ( .OUT(na773_1), .CLK(na2414_1), .EN(na154_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na773_1_i) );
// C_AND/D///      x116y38     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a774_1 ( .OUT(na774_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2403_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a774_2 ( .OUT(na774_1), .CLK(na2414_1), .EN(na154_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na774_1_i) );
// C_AND/D///      x116y42     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a775_1 ( .OUT(na775_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a775_2 ( .OUT(na775_1), .CLK(na2414_1), .EN(na154_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na775_1_i) );
// C_///AND/D      x119y50     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a776_4 ( .OUT(na776_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a776_5 ( .OUT(na776_2), .CLK(na2414_1), .EN(na154_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na776_2_i) );
// C_AND/D///      x122y50     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a777_1 ( .OUT(na777_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a777_2 ( .OUT(na777_1), .CLK(na2414_1), .EN(na154_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na777_1_i) );
// C_///AND/D      x133y70     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a778_4 ( .OUT(na778_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a778_5 ( .OUT(na778_2), .CLK(na2414_1), .EN(na154_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na778_2_i) );
// C_///AND/D      x126y68     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a779_4 ( .OUT(na779_2_i), .IN1(na2408_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a779_5 ( .OUT(na779_2), .CLK(na2414_1), .EN(na154_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na779_2_i) );
// C_///AND/D      x111y71     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a780_4 ( .OUT(na780_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a780_5 ( .OUT(na780_2), .CLK(na2414_1), .EN(na154_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na780_2_i) );
// C_AND/D///      x123y73     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a781_1 ( .OUT(na781_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a781_2 ( .OUT(na781_1), .CLK(na2414_1), .EN(na154_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na781_1_i) );
// C_AND/D///      x116y32     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a782_1 ( .OUT(na782_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2401_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a782_2 ( .OUT(na782_1), .CLK(na2414_1), .EN(na155_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na782_1_i) );
// C_AND/D///      x120y35     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a783_1 ( .OUT(na783_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a783_2 ( .OUT(na783_1), .CLK(na2414_1), .EN(na155_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na783_1_i) );
// C_///AND/D      x119y45     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a784_4 ( .OUT(na784_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a784_5 ( .OUT(na784_2), .CLK(na2414_1), .EN(na155_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na784_2_i) );
// C_///AND/D      x119y43     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a785_4 ( .OUT(na785_2_i), .IN1(1'b1), .IN2(na2404_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a785_5 ( .OUT(na785_2), .CLK(na2414_1), .EN(na155_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na785_2_i) );
// C_///AND/D      x120y51     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a786_4 ( .OUT(na786_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a786_5 ( .OUT(na786_2), .CLK(na2414_1), .EN(na155_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na786_2_i) );
// C_AND/D///      x125y49     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a787_1 ( .OUT(na787_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a787_2 ( .OUT(na787_1), .CLK(na2414_1), .EN(na155_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na787_1_i) );
// C_///AND/D      x134y71     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a788_4 ( .OUT(na788_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a788_5 ( .OUT(na788_2), .CLK(na2414_1), .EN(na155_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na788_2_i) );
// C_AND/D///      x121y65     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a789_1 ( .OUT(na789_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a789_2 ( .OUT(na789_1), .CLK(na2414_1), .EN(na155_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na789_1_i) );
// C_AND/D///      x114y76     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a790_1 ( .OUT(na790_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2409_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a790_2 ( .OUT(na790_1), .CLK(na2414_1), .EN(na155_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na790_1_i) );
// C_AND/D///      x128y76     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a791_1 ( .OUT(na791_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a791_2 ( .OUT(na791_1), .CLK(na2414_1), .EN(na155_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na791_1_i) );
// C_///AND/D      x116y29     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a792_4 ( .OUT(na792_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a792_5 ( .OUT(na792_2), .CLK(na2414_1), .EN(na156_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na792_2_i) );
// C_///AND/D      x122y38     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a793_4 ( .OUT(na793_2_i), .IN1(na2402_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a793_5 ( .OUT(na793_2), .CLK(na2414_1), .EN(na156_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na793_2_i) );
// C_///AND/D      x117y50     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a794_4 ( .OUT(na794_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a794_5 ( .OUT(na794_2), .CLK(na2414_1), .EN(na156_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na794_2_i) );
// C_AND/D///      x117y42     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a795_1 ( .OUT(na795_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a795_2 ( .OUT(na795_1), .CLK(na2414_1), .EN(na156_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na795_1_i) );
// C_AND/D///      x114y50     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a796_1 ( .OUT(na796_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2405_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a796_2 ( .OUT(na796_1), .CLK(na2414_1), .EN(na156_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na796_1_i) );
// C_AND/D///      x125y50     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a797_1 ( .OUT(na797_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a797_2 ( .OUT(na797_1), .CLK(na2414_1), .EN(na156_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na797_1_i) );
// C_///AND/D      x134y74     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a798_4 ( .OUT(na798_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a798_5 ( .OUT(na798_2), .CLK(na2414_1), .EN(na156_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na798_2_i) );
// C_AND/D///      x121y68     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a799_1 ( .OUT(na799_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a799_2 ( .OUT(na799_1), .CLK(na2414_1), .EN(na156_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na799_1_i) );
// C_///AND/D      x114y71     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a800_4 ( .OUT(na800_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a800_5 ( .OUT(na800_2), .CLK(na2414_1), .EN(na156_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na800_2_i) );
// C_///AND/D      x124y77     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a801_4 ( .OUT(na801_2_i), .IN1(1'b1), .IN2(na2410_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a801_5 ( .OUT(na801_2), .CLK(na2414_1), .EN(na156_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na801_2_i) );
// C_///AND/D      x114y34     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a802_4 ( .OUT(na802_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a802_5 ( .OUT(na802_2), .CLK(na2414_1), .EN(na157_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na802_2_i) );
// C_AND/D///      x120y37     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a803_1 ( .OUT(na803_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a803_2 ( .OUT(na803_1), .CLK(na2414_1), .EN(na157_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na803_1_i) );
// C_AND/D///      x118y35     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a804_1 ( .OUT(na804_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2403_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a804_2 ( .OUT(na804_1), .CLK(na2414_1), .EN(na157_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na804_1_i) );
// C_AND/D///      x115y43     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a805_1 ( .OUT(na805_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a805_2 ( .OUT(na805_1), .CLK(na2414_1), .EN(na157_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na805_1_i) );
// C_///AND/D      x116y49     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a806_4 ( .OUT(na806_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a806_5 ( .OUT(na806_2), .CLK(na2414_1), .EN(na157_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na806_2_i) );
// C_///AND/D      x124y49     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a807_4 ( .OUT(na807_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2406_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a807_5 ( .OUT(na807_2), .CLK(na2414_1), .EN(na157_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na807_2_i) );
// C_///AND/D      x126y67     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a808_4 ( .OUT(na808_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a808_5 ( .OUT(na808_2), .CLK(na2414_1), .EN(na157_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na808_2_i) );
// C_AND/D///      x123y68     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a809_1 ( .OUT(na809_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a809_2 ( .OUT(na809_1), .CLK(na2414_1), .EN(na157_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na809_1_i) );
// C_///AND/D      x114y67     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a810_4 ( .OUT(na810_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a810_5 ( .OUT(na810_2), .CLK(na2414_1), .EN(na157_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na810_2_i) );
// C_AND/D///      x125y75     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a811_1 ( .OUT(na811_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a811_2 ( .OUT(na811_1), .CLK(na2414_1), .EN(na157_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na811_1_i) );
// C_AND/D///      x116y31     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a812_1 ( .OUT(na812_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2401_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a812_2 ( .OUT(na812_1), .CLK(na2414_1), .EN(na158_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na812_1_i) );
// C_AND/D///      x120y40     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a813_1 ( .OUT(na813_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a813_2 ( .OUT(na813_1), .CLK(na2414_1), .EN(na158_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na813_1_i) );
// C_///AND/D      x118y42     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a814_4 ( .OUT(na814_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a814_5 ( .OUT(na814_2), .CLK(na2414_1), .EN(na158_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na814_2_i) );
// C_///AND/D      x117y46     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a815_4 ( .OUT(na815_2_i), .IN1(1'b1), .IN2(na2404_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a815_5 ( .OUT(na815_2), .CLK(na2414_1), .EN(na158_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na815_2_i) );
// C_///AND/D      x118y54     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a816_4 ( .OUT(na816_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a816_5 ( .OUT(na816_2), .CLK(na2414_1), .EN(na158_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na816_2_i) );
// C_AND/D///      x126y52     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a817_1 ( .OUT(na817_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a817_2 ( .OUT(na817_1), .CLK(na2414_1), .EN(na158_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na817_1_i) );
// C_AND/D///      x126y64     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a818_1 ( .OUT(na818_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2407_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a818_2 ( .OUT(na818_1), .CLK(na2414_1), .EN(na158_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na818_1_i) );
// C_AND/D///      x123y69     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a819_1 ( .OUT(na819_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a819_2 ( .OUT(na819_1), .CLK(na2414_1), .EN(na158_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na819_1_i) );
// C_///AND/D      x112y70     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a820_4 ( .OUT(na820_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a820_5 ( .OUT(na820_2), .CLK(na2414_1), .EN(na158_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na820_2_i) );
// C_AND/D///      x129y76     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a821_1 ( .OUT(na821_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a821_2 ( .OUT(na821_1), .CLK(na2414_1), .EN(na158_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na821_1_i) );
// C_///AND/D      x117y30     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a822_4 ( .OUT(na822_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a822_5 ( .OUT(na822_2), .CLK(na2414_1), .EN(na159_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na822_2_i) );
// C_///AND/D      x121y41     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a823_4 ( .OUT(na823_2_i), .IN1(na2402_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a823_5 ( .OUT(na823_2), .CLK(na2414_1), .EN(na159_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na823_2_i) );
// C_///AND/D      x119y39     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a824_4 ( .OUT(na824_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a824_5 ( .OUT(na824_2), .CLK(na2414_1), .EN(na159_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na824_2_i) );
// C_AND/D///      x116y43     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a825_1 ( .OUT(na825_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a825_2 ( .OUT(na825_1), .CLK(na2414_1), .EN(na159_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na825_1_i) );
// C_AND/D///      x113y47     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a826_1 ( .OUT(na826_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2405_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a826_2 ( .OUT(na826_1), .CLK(na2414_1), .EN(na159_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na826_1_i) );
// C_AND/D///      x125y51     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a827_1 ( .OUT(na827_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a827_2 ( .OUT(na827_1), .CLK(na2414_1), .EN(na159_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na827_1_i) );
// C_///AND/D      x129y65     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a828_4 ( .OUT(na828_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a828_5 ( .OUT(na828_2), .CLK(na2414_1), .EN(na159_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na828_2_i) );
// C_///AND/D      x124y70     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a829_4 ( .OUT(na829_2_i), .IN1(na2408_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a829_5 ( .OUT(na829_2), .CLK(na2414_1), .EN(na159_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na829_2_i) );
// C_///AND/D      x109y71     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a830_4 ( .OUT(na830_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a830_5 ( .OUT(na830_2), .CLK(na2414_1), .EN(na159_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na830_2_i) );
// C_AND/D///      x128y73     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a831_1 ( .OUT(na831_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a831_2 ( .OUT(na831_1), .CLK(na2414_1), .EN(na159_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na831_1_i) );
// C_///AND/D      x119y31     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a832_4 ( .OUT(na832_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a832_5 ( .OUT(na832_2), .CLK(na2414_1), .EN(na160_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na832_2_i) );
// C_AND/D///      x119y40     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a833_1 ( .OUT(na833_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a833_2 ( .OUT(na833_1), .CLK(na2414_1), .EN(na160_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na833_1_i) );
// C_AND/D///      x119y36     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a834_1 ( .OUT(na834_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2403_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a834_2 ( .OUT(na834_1), .CLK(na2414_1), .EN(na160_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na834_1_i) );
// C_AND/D///      x118y44     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a835_1 ( .OUT(na835_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a835_2 ( .OUT(na835_1), .CLK(na2414_1), .EN(na160_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na835_1_i) );
// C_///AND/D      x113y52     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a836_4 ( .OUT(na836_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a836_5 ( .OUT(na836_2), .CLK(na2414_1), .EN(na160_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na836_2_i) );
// C_///AND/D      x119y52     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a837_4 ( .OUT(na837_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2406_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a837_5 ( .OUT(na837_2), .CLK(na2414_1), .EN(na160_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na837_2_i) );
// C_///AND/D      x131y66     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a838_4 ( .OUT(na838_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a838_5 ( .OUT(na838_2), .CLK(na2414_1), .EN(na160_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na838_2_i) );
// C_AND/D///      x128y69     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a839_1 ( .OUT(na839_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a839_2 ( .OUT(na839_1), .CLK(na2414_1), .EN(na160_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na839_1_i) );
// C_AND/D///      x111y76     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a840_1 ( .OUT(na840_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2409_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a840_2 ( .OUT(na840_1), .CLK(na2414_1), .EN(na160_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na840_1_i) );
// C_AND/D///      x130y76     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a841_1 ( .OUT(na841_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a841_2 ( .OUT(na841_1), .CLK(na2414_1), .EN(na160_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na841_1_i) );
// C_///AND/D      x123y32     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a842_4 ( .OUT(na842_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a842_5 ( .OUT(na842_2), .CLK(na2414_1), .EN(na161_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na842_2_i) );
// C_AND/D///      x119y47     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a843_1 ( .OUT(na843_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a843_2 ( .OUT(na843_1), .CLK(na2414_1), .EN(na161_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na843_1_i) );
// C_///AND/D      x120y41     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a844_4 ( .OUT(na844_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a844_5 ( .OUT(na844_2), .CLK(na2414_1), .EN(na161_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na844_2_i) );
// C_///AND/D      x122y45     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a845_4 ( .OUT(na845_2_i), .IN1(1'b1), .IN2(na2404_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a845_5 ( .OUT(na845_2), .CLK(na2414_1), .EN(na161_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na845_2_i) );
// C_///AND/D      x113y55     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a846_4 ( .OUT(na846_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a846_5 ( .OUT(na846_2), .CLK(na2414_1), .EN(na161_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na846_2_i) );
// C_AND/D///      x123y52     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a847_1 ( .OUT(na847_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a847_2 ( .OUT(na847_1), .CLK(na2414_1), .EN(na161_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na847_1_i) );
// C_AND/D///      x131y65     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a848_1 ( .OUT(na848_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2407_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a848_2 ( .OUT(na848_1), .CLK(na2414_1), .EN(na161_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na848_1_i) );
// C_AND/D///      x123y71     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a849_1 ( .OUT(na849_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a849_2 ( .OUT(na849_1), .CLK(na2414_1), .EN(na161_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na849_1_i) );
// C_///AND/D      x118y73     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a850_4 ( .OUT(na850_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a850_5 ( .OUT(na850_2), .CLK(na2414_1), .EN(na161_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na850_2_i) );
// C_///AND/D      x126y79     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a851_4 ( .OUT(na851_2_i), .IN1(1'b1), .IN2(na2410_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a851_5 ( .OUT(na851_2), .CLK(na2414_1), .EN(na161_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na851_2_i) );
// C_///AND/D      x119y34     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a852_4 ( .OUT(na852_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a852_5 ( .OUT(na852_2), .CLK(na2414_1), .EN(na151_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na852_2_i) );
// C_AND/D///      x121y35     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a853_1 ( .OUT(na853_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a853_2 ( .OUT(na853_1), .CLK(na2414_1), .EN(na151_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na853_1_i) );
// C_///AND/D      x118y45     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a854_4 ( .OUT(na854_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a854_5 ( .OUT(na854_2), .CLK(na2414_1), .EN(na151_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na854_2_i) );
// C_AND/D///      x118y43     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a855_1 ( .OUT(na855_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a855_2 ( .OUT(na855_1), .CLK(na2414_1), .EN(na151_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na855_1_i) );
// C_AND/D///      x113y51     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a856_1 ( .OUT(na856_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2405_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a856_2 ( .OUT(na856_1), .CLK(na2414_1), .EN(na151_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na856_1_i) );
// C_AND/D///      x128y51     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a857_1 ( .OUT(na857_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a857_2 ( .OUT(na857_1), .CLK(na2414_1), .EN(na151_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na857_1_i) );
// C_///AND/D      x133y71     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a858_4 ( .OUT(na858_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a858_5 ( .OUT(na858_2), .CLK(na2414_1), .EN(na151_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na858_2_i) );
// C_///AND/D      x124y67     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a859_4 ( .OUT(na859_2_i), .IN1(na2408_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a859_5 ( .OUT(na859_2), .CLK(na2414_1), .EN(na151_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na859_2_i) );
// C_///AND/D      x113y70     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a860_4 ( .OUT(na860_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a860_5 ( .OUT(na860_2), .CLK(na2414_1), .EN(na151_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na860_2_i) );
// C_AND/D///      x125y76     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a861_1 ( .OUT(na861_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a861_2 ( .OUT(na861_1), .CLK(na2414_1), .EN(na151_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na861_1_i) );
// C_AND/D///      x118y32     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a862_1 ( .OUT(na862_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2401_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a862_2 ( .OUT(na862_1), .CLK(na2414_1), .EN(na163_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na862_1_i) );
// C_AND/D///      x120y43     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a863_1 ( .OUT(na863_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a863_2 ( .OUT(na863_1), .CLK(na2414_1), .EN(na163_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na863_1_i) );
// C_///AND/D      x121y45     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a864_4 ( .OUT(na864_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a864_5 ( .OUT(na864_2), .CLK(na2414_1), .EN(na163_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na864_2_i) );
// C_AND/D///      x119y41     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a865_1 ( .OUT(na865_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a865_2 ( .OUT(na865_1), .CLK(na2414_1), .EN(na163_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na865_1_i) );
// C_///AND/D      x114y55     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a866_4 ( .OUT(na866_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a866_5 ( .OUT(na866_2), .CLK(na2414_1), .EN(na163_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na866_2_i) );
// C_///AND/D      x124y50     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a867_4 ( .OUT(na867_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2406_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a867_5 ( .OUT(na867_2), .CLK(na2414_1), .EN(na163_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na867_2_i) );
// C_///AND/D      x138y71     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a868_4 ( .OUT(na868_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a868_5 ( .OUT(na868_2), .CLK(na2414_1), .EN(na163_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na868_2_i) );
// C_AND/D///      x126y71     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a869_1 ( .OUT(na869_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a869_2 ( .OUT(na869_1), .CLK(na2414_1), .EN(na163_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na869_1_i) );
// C_AND/D///      x115y75     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a870_1 ( .OUT(na870_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2409_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a870_2 ( .OUT(na870_1), .CLK(na2414_1), .EN(na163_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na870_1_i) );
// C_AND/D///      x125y77     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a871_1 ( .OUT(na871_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a871_2 ( .OUT(na871_1), .CLK(na2414_1), .EN(na163_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na871_1_i) );
// C_///AND/D      x118y33     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a872_4 ( .OUT(na872_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a872_5 ( .OUT(na872_2), .CLK(na2414_1), .EN(na164_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na872_2_i) );
// C_///AND/D      x122y42     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a873_4 ( .OUT(na873_2_i), .IN1(na2402_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a873_5 ( .OUT(na873_2), .CLK(na2414_1), .EN(na164_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na873_2_i) );
// C_///AND/D      x121y48     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a874_4 ( .OUT(na874_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a874_5 ( .OUT(na874_2), .CLK(na2414_1), .EN(na164_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na874_2_i) );
// C_AND/D///      x119y42     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a875_1 ( .OUT(na875_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a875_2 ( .OUT(na875_1), .CLK(na2414_1), .EN(na164_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na875_1_i) );
// C_///AND/D      x116y58     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a876_4 ( .OUT(na876_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a876_5 ( .OUT(na876_2), .CLK(na2414_1), .EN(na164_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na876_2_i) );
// C_AND/D///      x124y51     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a877_1 ( .OUT(na877_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a877_2 ( .OUT(na877_1), .CLK(na2414_1), .EN(na164_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na877_1_i) );
// C_AND/D///      x132y66     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a878_1 ( .OUT(na878_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2407_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a878_2 ( .OUT(na878_1), .CLK(na2414_1), .EN(na164_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na878_1_i) );
// C_AND/D///      x124y72     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a879_1 ( .OUT(na879_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a879_2 ( .OUT(na879_1), .CLK(na2414_1), .EN(na164_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na879_1_i) );
// C_///AND/D      x123y74     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a880_4 ( .OUT(na880_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a880_5 ( .OUT(na880_2), .CLK(na2414_1), .EN(na164_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na880_2_i) );
// C_///AND/D      x123y82     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a881_4 ( .OUT(na881_2_i), .IN1(1'b1), .IN2(na2410_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a881_5 ( .OUT(na881_2), .CLK(na2414_1), .EN(na164_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na881_2_i) );
// C_///AND/D      x122y34     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a882_4 ( .OUT(na882_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a882_5 ( .OUT(na882_2), .CLK(na2414_1), .EN(na165_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na882_2_i) );
// C_AND/D///      x123y41     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a883_1 ( .OUT(na883_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a883_2 ( .OUT(na883_1), .CLK(na2414_1), .EN(na165_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na883_1_i) );
// C_AND/D///      x115y36     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a884_1 ( .OUT(na884_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2403_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a884_2 ( .OUT(na884_1), .CLK(na2414_1), .EN(na165_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na884_1_i) );
// C_AND/D///      x121y43     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a885_1 ( .OUT(na885_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a885_2 ( .OUT(na885_1), .CLK(na2414_1), .EN(na165_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na885_1_i) );
// C_///AND/D      x119y54     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a886_4 ( .OUT(na886_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a886_5 ( .OUT(na886_2), .CLK(na2414_1), .EN(na165_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na886_2_i) );
// C_AND/D///      x129y54     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a887_1 ( .OUT(na887_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a887_2 ( .OUT(na887_1), .CLK(na2414_1), .EN(na165_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na887_1_i) );
// C_///AND/D      x134y65     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a888_4 ( .OUT(na888_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a888_5 ( .OUT(na888_2), .CLK(na2414_1), .EN(na165_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na888_2_i) );
// C_///AND/D      x123y76     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a889_4 ( .OUT(na889_2_i), .IN1(na2408_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a889_5 ( .OUT(na889_2), .CLK(na2414_1), .EN(na165_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na889_2_i) );
// C_///AND/D      x113y77     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a890_4 ( .OUT(na890_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a890_5 ( .OUT(na890_2), .CLK(na2414_1), .EN(na165_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na890_2_i) );
// C_AND/D///      x124y78     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a891_1 ( .OUT(na891_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a891_2 ( .OUT(na891_1), .CLK(na2414_1), .EN(na165_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na891_1_i) );
// C_AND/D///      x120y31     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a892_1 ( .OUT(na892_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2401_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a892_2 ( .OUT(na892_1), .CLK(na2414_1), .EN(na166_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na892_1_i) );
// C_AND/D///      x121y42     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a893_1 ( .OUT(na893_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a893_2 ( .OUT(na893_1), .CLK(na2414_1), .EN(na166_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na893_1_i) );
// C_///AND/D      x117y41     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a894_4 ( .OUT(na894_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a894_5 ( .OUT(na894_2), .CLK(na2414_1), .EN(na166_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na894_2_i) );
// C_///AND/D      x121y44     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a895_4 ( .OUT(na895_2_i), .IN1(1'b1), .IN2(na2404_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a895_5 ( .OUT(na895_2), .CLK(na2414_1), .EN(na166_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na895_2_i) );
// C_///AND/D      x119y53     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a896_4 ( .OUT(na896_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a896_5 ( .OUT(na896_2), .CLK(na2414_1), .EN(na166_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na896_2_i) );
// C_AND/D///      x131y53     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a897_1 ( .OUT(na897_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a897_2 ( .OUT(na897_1), .CLK(na2414_1), .EN(na166_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na897_1_i) );
// C_///AND/D      x136y72     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a898_4 ( .OUT(na898_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a898_5 ( .OUT(na898_2), .CLK(na2414_1), .EN(na166_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na898_2_i) );
// C_AND/D///      x121y71     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a899_1 ( .OUT(na899_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a899_2 ( .OUT(na899_1), .CLK(na2414_1), .EN(na166_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na899_1_i) );
// C_AND/D///      x113y82     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a900_1 ( .OUT(na900_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2409_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a900_2 ( .OUT(na900_1), .CLK(na2414_1), .EN(na166_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na900_1_i) );
// C_AND/D///      x126y77     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a901_1 ( .OUT(na901_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a901_2 ( .OUT(na901_1), .CLK(na2414_1), .EN(na166_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na901_1_i) );
// C_///AND/D      x121y36     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a902_4 ( .OUT(na902_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a902_5 ( .OUT(na902_2), .CLK(na2414_1), .EN(na167_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na902_2_i) );
// C_///AND/D      x122y43     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a903_4 ( .OUT(na903_2_i), .IN1(na2402_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a903_5 ( .OUT(na903_2), .CLK(na2414_1), .EN(na167_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na903_2_i) );
// C_///AND/D      x116y44     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a904_4 ( .OUT(na904_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a904_5 ( .OUT(na904_2), .CLK(na2414_1), .EN(na167_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na904_2_i) );
// C_AND/D///      x120y45     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a905_1 ( .OUT(na905_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a905_2 ( .OUT(na905_1), .CLK(na2414_1), .EN(na167_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na905_1_i) );
// C_AND/D///      x114y54     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a906_1 ( .OUT(na906_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2405_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a906_2 ( .OUT(na906_1), .CLK(na2414_1), .EN(na167_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na906_1_i) );
// C_AND/D///      x128y54     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a907_1 ( .OUT(na907_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a907_2 ( .OUT(na907_1), .CLK(na2414_1), .EN(na167_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na907_1_i) );
// C_///AND/D      x137y69     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a908_4 ( .OUT(na908_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a908_5 ( .OUT(na908_2), .CLK(na2414_1), .EN(na167_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na908_2_i) );
// C_AND/D///      x122y72     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a909_1 ( .OUT(na909_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a909_2 ( .OUT(na909_1), .CLK(na2414_1), .EN(na167_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na909_1_i) );
// C_///AND/D      x118y81     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a910_4 ( .OUT(na910_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a910_5 ( .OUT(na910_2), .CLK(na2414_1), .EN(na167_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na910_2_i) );
// C_///AND/D      x127y80     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a911_4 ( .OUT(na911_2_i), .IN1(1'b1), .IN2(na2410_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a911_5 ( .OUT(na911_2), .CLK(na2414_1), .EN(na167_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na911_2_i) );
// C_///AND/D      x119y35     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a912_4 ( .OUT(na912_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a912_5 ( .OUT(na912_2), .CLK(na2414_1), .EN(na162_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na912_2_i) );
// C_AND/D///      x123y44     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a913_1 ( .OUT(na913_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a913_2 ( .OUT(na913_1), .CLK(na2414_1), .EN(na162_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na913_1_i) );
// C_AND/D///      x118y38     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a914_1 ( .OUT(na914_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2403_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a914_2 ( .OUT(na914_1), .CLK(na2414_1), .EN(na162_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na914_1_i) );
// C_AND/D///      x120y42     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a915_1 ( .OUT(na915_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a915_2 ( .OUT(na915_1), .CLK(na2414_1), .EN(na162_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na915_1_i) );
// C_///AND/D      x113y54     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a916_4 ( .OUT(na916_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a916_5 ( .OUT(na916_2), .CLK(na2414_1), .EN(na162_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na916_2_i) );
// C_///AND/D      x121y53     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a917_4 ( .OUT(na917_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2406_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a917_5 ( .OUT(na917_2), .CLK(na2414_1), .EN(na162_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na917_2_i) );
// C_///AND/D      x137y74     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a918_4 ( .OUT(na918_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a918_5 ( .OUT(na918_2), .CLK(na2414_1), .EN(na162_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na918_2_i) );
// C_AND/D///      x125y72     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a919_1 ( .OUT(na919_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a919_2 ( .OUT(na919_1), .CLK(na2414_1), .EN(na162_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na919_1_i) );
// C_///AND/D      x122y78     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a920_4 ( .OUT(na920_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a920_5 ( .OUT(na920_2), .CLK(na2414_1), .EN(na162_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na920_2_i) );
// C_AND/D///      x122y78     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a921_1 ( .OUT(na921_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a921_2 ( .OUT(na921_1), .CLK(na2414_1), .EN(na162_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na921_1_i) );
// C_AND/D///      x127y31     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a922_1 ( .OUT(na922_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2401_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a922_2 ( .OUT(na922_1), .CLK(na2414_1), .EN(na186_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na922_1_i) );
// C_AND/D///      x126y36     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a923_1 ( .OUT(na923_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a923_2 ( .OUT(na923_1), .CLK(na2414_1), .EN(na186_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na923_1_i) );
// C_///AND/D      x114y43     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a924_4 ( .OUT(na924_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a924_5 ( .OUT(na924_2), .CLK(na2414_1), .EN(na186_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na924_2_i) );
// C_///AND/D      x122y47     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a925_4 ( .OUT(na925_2_i), .IN1(1'b1), .IN2(na2404_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a925_5 ( .OUT(na925_2), .CLK(na2414_1), .EN(na186_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na925_2_i) );
// C_///AND/D      x122y51     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a926_4 ( .OUT(na926_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a926_5 ( .OUT(na926_2), .CLK(na2414_1), .EN(na186_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na926_2_i) );
// C_AND/D///      x115y57     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a927_1 ( .OUT(na927_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a927_2 ( .OUT(na927_1), .CLK(na2414_1), .EN(na186_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na927_1_i) );
// C_AND/D///      x116y63     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a928_1 ( .OUT(na928_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2407_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a928_2 ( .OUT(na928_1), .CLK(na2414_1), .EN(na186_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na928_1_i) );
// C_AND/D///      x113y68     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a929_1 ( .OUT(na929_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a929_2 ( .OUT(na929_1), .CLK(na2414_1), .EN(na186_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na929_1_i) );
// C_///AND/D      x124y82     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a930_4 ( .OUT(na930_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a930_5 ( .OUT(na930_2), .CLK(na2414_1), .EN(na186_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na930_2_i) );
// C_AND/D///      x140y69     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a931_1 ( .OUT(na931_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a931_2 ( .OUT(na931_1), .CLK(na2414_1), .EN(na186_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na931_1_i) );
// C_///AND/D      x123y31     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a932_4 ( .OUT(na932_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a932_5 ( .OUT(na932_2), .CLK(na2414_1), .EN(na172_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na932_2_i) );
// C_///AND/D      x121y34     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a933_4 ( .OUT(na933_2_i), .IN1(na2402_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a933_5 ( .OUT(na933_2), .CLK(na2414_1), .EN(na172_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na933_2_i) );
// C_///AND/D      x114y47     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a934_4 ( .OUT(na934_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a934_5 ( .OUT(na934_2), .CLK(na2414_1), .EN(na172_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na934_2_i) );
// C_AND/D///      x112y45     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a935_1 ( .OUT(na935_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a935_2 ( .OUT(na935_1), .CLK(na2414_1), .EN(na172_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na935_1_i) );
// C_AND/D///      x111y53     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a936_1 ( .OUT(na936_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2405_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a936_2 ( .OUT(na936_1), .CLK(na2414_1), .EN(na172_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na936_1_i) );
// C_AND/D///      x115y55     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a937_1 ( .OUT(na937_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a937_2 ( .OUT(na937_1), .CLK(na2414_1), .EN(na172_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na937_1_i) );
// C_///AND/D      x117y67     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a938_4 ( .OUT(na938_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a938_5 ( .OUT(na938_2), .CLK(na2414_1), .EN(na172_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na938_2_i) );
// C_///AND/D      x114y65     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a939_4 ( .OUT(na939_2_i), .IN1(na2408_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a939_5 ( .OUT(na939_2), .CLK(na2414_1), .EN(na172_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na939_2_i) );
// C_///AND/D      x119y75     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a940_4 ( .OUT(na940_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a940_5 ( .OUT(na940_2), .CLK(na2414_1), .EN(na172_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na940_2_i) );
// C_AND/D///      x135y74     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a941_1 ( .OUT(na941_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a941_2 ( .OUT(na941_1), .CLK(na2414_1), .EN(na172_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na941_1_i) );
// C_///AND/D      x126y30     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a942_4 ( .OUT(na942_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a942_5 ( .OUT(na942_2), .CLK(na2414_1), .EN(na173_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na942_2_i) );
// C_AND/D///      x120y33     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a943_1 ( .OUT(na943_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a943_2 ( .OUT(na943_1), .CLK(na2414_1), .EN(na173_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na943_1_i) );
// C_AND/D///      x111y40     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a944_1 ( .OUT(na944_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2403_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a944_2 ( .OUT(na944_1), .CLK(na2414_1), .EN(na173_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na944_1_i) );
// C_AND/D///      x115y46     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a945_1 ( .OUT(na945_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a945_2 ( .OUT(na945_1), .CLK(na2414_1), .EN(na173_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na945_1_i) );
// C_///AND/D      x118y50     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a946_4 ( .OUT(na946_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a946_5 ( .OUT(na946_2), .CLK(na2414_1), .EN(na173_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na946_2_i) );
// C_///AND/D      x122y56     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a947_4 ( .OUT(na947_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2406_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a947_5 ( .OUT(na947_2), .CLK(na2414_1), .EN(na173_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na947_2_i) );
// C_///AND/D      x116y70     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a948_4 ( .OUT(na948_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a948_5 ( .OUT(na948_2), .CLK(na2414_1), .EN(na173_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na948_2_i) );
// C_AND/D///      x111y66     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a949_1 ( .OUT(na949_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a949_2 ( .OUT(na949_1), .CLK(na2414_1), .EN(na173_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na949_1_i) );
// C_AND/D///      x116y78     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a950_1 ( .OUT(na950_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2409_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a950_2 ( .OUT(na950_1), .CLK(na2414_1), .EN(na173_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na950_1_i) );
// C_AND/D///      x136y75     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a951_1 ( .OUT(na951_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a951_2 ( .OUT(na951_1), .CLK(na2414_1), .EN(na173_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na951_1_i) );
// C_///AND/D      x126y31     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a952_4 ( .OUT(na952_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a952_5 ( .OUT(na952_2), .CLK(na2414_1), .EN(na174_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na952_2_i) );
// C_AND/D///      x124y34     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a953_1 ( .OUT(na953_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a953_2 ( .OUT(na953_1), .CLK(na2414_1), .EN(na174_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na953_1_i) );
// C_///AND/D      x117y47     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a954_4 ( .OUT(na954_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a954_5 ( .OUT(na954_2), .CLK(na2414_1), .EN(na174_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na954_2_i) );
// C_///AND/D      x121y49     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a955_4 ( .OUT(na955_2_i), .IN1(1'b1), .IN2(na2404_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a955_5 ( .OUT(na955_2), .CLK(na2414_1), .EN(na174_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na955_2_i) );
// C_///AND/D      x116y45     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a956_4 ( .OUT(na956_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a956_5 ( .OUT(na956_2), .CLK(na2414_1), .EN(na174_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na956_2_i) );
// C_AND/D///      x112y55     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a957_1 ( .OUT(na957_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a957_2 ( .OUT(na957_1), .CLK(na2414_1), .EN(na174_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na957_1_i) );
// C_AND/D///      x118y65     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a958_1 ( .OUT(na958_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2407_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a958_2 ( .OUT(na958_1), .CLK(na2414_1), .EN(na174_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na958_1_i) );
// C_AND/D///      x109y65     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a959_1 ( .OUT(na959_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a959_2 ( .OUT(na959_1), .CLK(na2414_1), .EN(na174_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na959_1_i) );
// C_///AND/D      x122y79     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a960_4 ( .OUT(na960_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a960_5 ( .OUT(na960_2), .CLK(na2414_1), .EN(na174_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na960_2_i) );
// C_///AND/D      x136y76     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a961_4 ( .OUT(na961_2_i), .IN1(1'b1), .IN2(na2410_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a961_5 ( .OUT(na961_2), .CLK(na2414_1), .EN(na174_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na961_2_i) );
// C_///AND/D      x132y32     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a962_4 ( .OUT(na962_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a962_5 ( .OUT(na962_2), .CLK(na2414_1), .EN(na175_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na962_2_i) );
// C_AND/D///      x124y36     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a963_1 ( .OUT(na963_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a963_2 ( .OUT(na963_1), .CLK(na2414_1), .EN(na175_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na963_1_i) );
// C_///AND/D      x115y47     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a964_4 ( .OUT(na964_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a964_5 ( .OUT(na964_2), .CLK(na2414_1), .EN(na175_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na964_2_i) );
// C_AND/D///      x116y47     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a965_1 ( .OUT(na965_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a965_2 ( .OUT(na965_1), .CLK(na2414_1), .EN(na175_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na965_1_i) );
// C_AND/D///      x114y53     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a966_1 ( .OUT(na966_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2405_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a966_2 ( .OUT(na966_1), .CLK(na2414_1), .EN(na175_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na966_1_i) );
// C_AND/D///      x116y52     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a967_1 ( .OUT(na967_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a967_2 ( .OUT(na967_1), .CLK(na2414_1), .EN(na175_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na967_1_i) );
// C_///AND/D      x122y64     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a968_4 ( .OUT(na968_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a968_5 ( .OUT(na968_2), .CLK(na2414_1), .EN(na175_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na968_2_i) );
// C_///AND/D      x113y67     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a969_4 ( .OUT(na969_2_i), .IN1(na2408_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a969_5 ( .OUT(na969_2), .CLK(na2414_1), .EN(na175_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na969_2_i) );
// C_///AND/D      x118y75     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a970_4 ( .OUT(na970_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a970_5 ( .OUT(na970_2), .CLK(na2414_1), .EN(na175_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na970_2_i) );
// C_AND/D///      x135y69     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a971_1 ( .OUT(na971_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a971_2 ( .OUT(na971_1), .CLK(na2414_1), .EN(na175_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na971_1_i) );
// C_AND/D///      x124y31     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a972_1 ( .OUT(na972_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2401_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a972_2 ( .OUT(na972_1), .CLK(na2414_1), .EN(na176_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na972_1_i) );
// C_AND/D///      x122y33     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a973_1 ( .OUT(na973_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a973_2 ( .OUT(na973_1), .CLK(na2414_1), .EN(na176_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na973_1_i) );
// C_///AND/D      x113y46     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a974_4 ( .OUT(na974_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a974_5 ( .OUT(na974_2), .CLK(na2414_1), .EN(na176_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na974_2_i) );
// C_AND/D///      x118y48     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a975_1 ( .OUT(na975_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a975_2 ( .OUT(na975_1), .CLK(na2414_1), .EN(na176_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na975_1_i) );
// C_///AND/D      x118y56     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a976_4 ( .OUT(na976_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a976_5 ( .OUT(na976_2), .CLK(na2414_1), .EN(na176_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na976_2_i) );
// C_///AND/D      x118y55     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a977_4 ( .OUT(na977_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2406_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a977_5 ( .OUT(na977_2), .CLK(na2414_1), .EN(na176_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na977_2_i) );
// C_///AND/D      x122y65     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a978_4 ( .OUT(na978_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a978_5 ( .OUT(na978_2), .CLK(na2414_1), .EN(na176_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na978_2_i) );
// C_AND/D///      x115y72     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a979_1 ( .OUT(na979_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a979_2 ( .OUT(na979_1), .CLK(na2414_1), .EN(na176_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na979_1_i) );
// C_AND/D///      x114y80     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a980_1 ( .OUT(na980_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2409_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a980_2 ( .OUT(na980_1), .CLK(na2414_1), .EN(na176_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na980_1_i) );
// C_AND/D///      x139y70     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a981_1 ( .OUT(na981_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a981_2 ( .OUT(na981_1), .CLK(na2414_1), .EN(na176_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na981_1_i) );
// C_///AND/D      x135y30     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a982_4 ( .OUT(na982_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a982_5 ( .OUT(na982_2), .CLK(na2414_1), .EN(na177_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na982_2_i) );
// C_///AND/D      x123y34     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a983_4 ( .OUT(na983_2_i), .IN1(na2402_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a983_5 ( .OUT(na983_2), .CLK(na2414_1), .EN(na177_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na983_2_i) );
// C_///AND/D      x112y49     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a984_4 ( .OUT(na984_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a984_5 ( .OUT(na984_2), .CLK(na2414_1), .EN(na177_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na984_2_i) );
// C_AND/D///      x115y49     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a985_1 ( .OUT(na985_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a985_2 ( .OUT(na985_1), .CLK(na2414_1), .EN(na177_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na985_1_i) );
// C_AND/D///      x113y57     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a986_1 ( .OUT(na986_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2405_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a986_2 ( .OUT(na986_1), .CLK(na2414_1), .EN(na177_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na986_1_i) );
// C_AND/D///      x115y50     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a987_1 ( .OUT(na987_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a987_2 ( .OUT(na987_1), .CLK(na2414_1), .EN(na177_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na987_1_i) );
// C_///AND/D      x119y68     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a988_4 ( .OUT(na988_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a988_5 ( .OUT(na988_2), .CLK(na2414_1), .EN(na177_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na988_2_i) );
// C_AND/D///      x116y71     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a989_1 ( .OUT(na989_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a989_2 ( .OUT(na989_1), .CLK(na2414_1), .EN(na177_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na989_1_i) );
// C_///AND/D      x119y77     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a990_4 ( .OUT(na990_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a990_5 ( .OUT(na990_2), .CLK(na2414_1), .EN(na177_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na990_2_i) );
// C_AND/D///      x140y71     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a991_1 ( .OUT(na991_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a991_2 ( .OUT(na991_1), .CLK(na2414_1), .EN(na177_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na991_1_i) );
// C_///AND/D      x133y31     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a992_4 ( .OUT(na992_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a992_5 ( .OUT(na992_2), .CLK(na2414_1), .EN(na178_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na992_2_i) );
// C_///AND/D      x123y35     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a993_4 ( .OUT(na993_2_i), .IN1(na2402_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a993_5 ( .OUT(na993_2), .CLK(na2414_1), .EN(na178_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na993_2_i) );
// C_///AND/D      x112y46     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a994_4 ( .OUT(na994_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a994_5 ( .OUT(na994_2), .CLK(na2414_1), .EN(na178_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na994_2_i) );
// C_AND/D///      x113y50     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a995_1 ( .OUT(na995_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a995_2 ( .OUT(na995_1), .CLK(na2414_1), .EN(na178_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na995_1_i) );
// C_///AND/D      x117y56     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a996_4 ( .OUT(na996_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a996_5 ( .OUT(na996_2), .CLK(na2414_1), .EN(na178_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na996_2_i) );
// C_AND/D///      x117y51     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a997_1 ( .OUT(na997_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a997_2 ( .OUT(na997_1), .CLK(na2414_1), .EN(na178_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na997_1_i) );
// C_///AND/D      x123y67     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a998_4 ( .OUT(na998_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a998_5 ( .OUT(na998_2), .CLK(na2414_1), .EN(na178_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na998_2_i) );
// C_AND/D///      x114y72     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a999_1 ( .OUT(na999_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a999_2 ( .OUT(na999_1), .CLK(na2414_1), .EN(na178_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na999_1_i) );
// C_AND/D///      x115y80     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1000_1 ( .OUT(na1000_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2409_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1000_2 ( .OUT(na1000_1), .CLK(na2414_1), .EN(na178_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1000_1_i) );
// C_AND/D///      x138y72     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1001_1 ( .OUT(na1001_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1001_2 ( .OUT(na1001_1), .CLK(na2414_1), .EN(na178_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1001_1_i) );
// C_///AND/D      x141y31     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1002_4 ( .OUT(na1002_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1002_5 ( .OUT(na1002_2), .CLK(na2414_1), .EN(na179_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1002_2_i) );
// C_AND/D///      x123y37     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1003_1 ( .OUT(na1003_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1003_2 ( .OUT(na1003_1), .CLK(na2414_1), .EN(na179_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1003_1_i) );
// C_///AND/D      x112y42     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1004_4 ( .OUT(na1004_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1004_5 ( .OUT(na1004_2), .CLK(na2414_1), .EN(na179_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1004_2_i) );
// C_AND/D///      x118y47     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1005_1 ( .OUT(na1005_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1005_2 ( .OUT(na1005_1), .CLK(na2414_1), .EN(na179_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1005_1_i) );
// C_///AND/D      x115y59     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1006_4 ( .OUT(na1006_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1006_5 ( .OUT(na1006_2), .CLK(na2414_1), .EN(na179_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1006_2_i) );
// C_///AND/D      x121y57     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1007_4 ( .OUT(na1007_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2406_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1007_5 ( .OUT(na1007_2), .CLK(na2414_1), .EN(na179_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1007_2_i) );
// C_///AND/D      x117y70     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1008_4 ( .OUT(na1008_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1008_5 ( .OUT(na1008_2), .CLK(na2414_1), .EN(na179_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1008_2_i) );
// C_AND/D///      x113y69     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1009_1 ( .OUT(na1009_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1009_2 ( .OUT(na1009_1), .CLK(na2414_1), .EN(na179_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1009_1_i) );
// C_///AND/D      x113y69     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1010_4 ( .OUT(na1010_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1010_5 ( .OUT(na1010_2), .CLK(na2414_1), .EN(na179_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1010_2_i) );
// C_AND/D///      x135y72     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1011_1 ( .OUT(na1011_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1011_2 ( .OUT(na1011_1), .CLK(na2414_1), .EN(na179_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1011_1_i) );
// C_///AND/D      x129y34     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1012_4 ( .OUT(na1012_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1012_5 ( .OUT(na1012_2), .CLK(na2414_1), .EN(na169_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1012_2_i) );
// C_AND/D///      x121y33     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1013_1 ( .OUT(na1013_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1013_2 ( .OUT(na1013_1), .CLK(na2414_1), .EN(na169_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1013_1_i) );
// C_AND/D///      x112y40     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1014_1 ( .OUT(na1014_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2403_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1014_2 ( .OUT(na1014_1), .CLK(na2414_1), .EN(na169_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1014_1_i) );
// C_AND/D///      x114y48     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1015_1 ( .OUT(na1015_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1015_2 ( .OUT(na1015_1), .CLK(na2414_1), .EN(na169_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1015_1_i) );
// C_///AND/D      x117y52     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1016_4 ( .OUT(na1016_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1016_5 ( .OUT(na1016_2), .CLK(na2414_1), .EN(na169_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1016_2_i) );
// C_AND/D///      x115y56     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1017_1 ( .OUT(na1017_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1017_2 ( .OUT(na1017_1), .CLK(na2414_1), .EN(na169_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1017_1_i) );
// C_///AND/D      x117y68     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1018_4 ( .OUT(na1018_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1018_5 ( .OUT(na1018_2), .CLK(na2414_1), .EN(na169_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1018_2_i) );
// C_AND/D///      x112y68     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1019_1 ( .OUT(na1019_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1019_2 ( .OUT(na1019_1), .CLK(na2414_1), .EN(na169_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1019_1_i) );
// C_///AND/D      x117y76     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1020_4 ( .OUT(na1020_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1020_5 ( .OUT(na1020_2), .CLK(na2414_1), .EN(na169_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1020_2_i) );
// C_///AND/D      x137y77     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1021_4 ( .OUT(na1021_2_i), .IN1(1'b1), .IN2(na2410_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1021_5 ( .OUT(na1021_2), .CLK(na2414_1), .EN(na169_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1021_2_i) );
// C_///AND/D      x142y33     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1022_4 ( .OUT(na1022_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1022_5 ( .OUT(na1022_2), .CLK(na2414_1), .EN(na181_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1022_2_i) );
// C_AND/D///      x122y37     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1023_1 ( .OUT(na1023_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1023_2 ( .OUT(na1023_1), .CLK(na2414_1), .EN(na181_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1023_1_i) );
// C_///AND/D      x111y44     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1024_4 ( .OUT(na1024_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1024_5 ( .OUT(na1024_2), .CLK(na2414_1), .EN(na181_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1024_2_i) );
// C_AND/D///      x117y45     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1025_1 ( .OUT(na1025_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1025_2 ( .OUT(na1025_1), .CLK(na2414_1), .EN(na181_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1025_1_i) );
// C_///AND/D      x118y57     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1026_4 ( .OUT(na1026_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1026_5 ( .OUT(na1026_2), .CLK(na2414_1), .EN(na181_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1026_2_i) );
// C_AND/D///      x120y55     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1027_1 ( .OUT(na1027_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1027_2 ( .OUT(na1027_1), .CLK(na2414_1), .EN(na181_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1027_1_i) );
// C_AND/D///      x116y66     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1028_1 ( .OUT(na1028_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2407_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1028_2 ( .OUT(na1028_1), .CLK(na2414_1), .EN(na181_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1028_1_i) );
// C_AND/D///      x112y69     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1029_1 ( .OUT(na1029_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1029_2 ( .OUT(na1029_1), .CLK(na2414_1), .EN(na181_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1029_1_i) );
// C_///AND/D      x116y67     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1030_4 ( .OUT(na1030_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1030_5 ( .OUT(na1030_2), .CLK(na2414_1), .EN(na181_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1030_2_i) );
// C_AND/D///      x136y70     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1031_1 ( .OUT(na1031_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1031_2 ( .OUT(na1031_1), .CLK(na2414_1), .EN(na181_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1031_1_i) );
// C_///AND/D      x142y32     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1032_4 ( .OUT(na1032_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1032_5 ( .OUT(na1032_2), .CLK(na2414_1), .EN(na182_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1032_2_i) );
// C_AND/D///      x122y40     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1033_1 ( .OUT(na1033_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1033_2 ( .OUT(na1033_1), .CLK(na2414_1), .EN(na182_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1033_1_i) );
// C_///AND/D      x109y43     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1034_4 ( .OUT(na1034_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1034_5 ( .OUT(na1034_2), .CLK(na2414_1), .EN(na182_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1034_2_i) );
// C_///AND/D      x121y50     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1035_4 ( .OUT(na1035_2_i), .IN1(1'b1), .IN2(na2404_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1035_5 ( .OUT(na1035_2), .CLK(na2414_1), .EN(na182_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1035_2_i) );
// C_///AND/D      x118y60     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1036_4 ( .OUT(na1036_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1036_5 ( .OUT(na1036_2), .CLK(na2414_1), .EN(na182_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1036_2_i) );
// C_AND/D///      x120y56     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1037_1 ( .OUT(na1037_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1037_2 ( .OUT(na1037_1), .CLK(na2414_1), .EN(na182_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1037_1_i) );
// C_///AND/D      x122y71     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1038_4 ( .OUT(na1038_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1038_5 ( .OUT(na1038_2), .CLK(na2414_1), .EN(na182_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1038_2_i) );
// C_AND/D///      x110y72     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1039_1 ( .OUT(na1039_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1039_2 ( .OUT(na1039_1), .CLK(na2414_1), .EN(na182_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1039_1_i) );
// C_///AND/D      x114y70     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1040_4 ( .OUT(na1040_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1040_5 ( .OUT(na1040_2), .CLK(na2414_1), .EN(na182_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1040_2_i) );
// C_AND/D///      x136y71     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1041_1 ( .OUT(na1041_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1041_2 ( .OUT(na1041_1), .CLK(na2414_1), .EN(na182_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1041_1_i) );
// C_AND/D///      x126y32     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1042_1 ( .OUT(na1042_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2401_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1042_2 ( .OUT(na1042_1), .CLK(na2414_1), .EN(na183_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1042_1_i) );
// C_AND/D///      x125y37     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1043_1 ( .OUT(na1043_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1043_2 ( .OUT(na1043_1), .CLK(na2414_1), .EN(na183_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1043_1_i) );
// C_///AND/D      x113y48     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1044_4 ( .OUT(na1044_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1044_5 ( .OUT(na1044_2), .CLK(na2414_1), .EN(na183_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1044_2_i) );
// C_AND/D///      x117y48     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1045_1 ( .OUT(na1045_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1045_2 ( .OUT(na1045_1), .CLK(na2414_1), .EN(na183_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1045_1_i) );
// C_///AND/D      x121y52     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1046_4 ( .OUT(na1046_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1046_5 ( .OUT(na1046_2), .CLK(na2414_1), .EN(na183_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1046_2_i) );
// C_AND/D///      x120y58     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1047_1 ( .OUT(na1047_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1047_2 ( .OUT(na1047_1), .CLK(na2414_1), .EN(na183_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1047_1_i) );
// C_///AND/D      x115y66     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1048_4 ( .OUT(na1048_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1048_5 ( .OUT(na1048_2), .CLK(na2414_1), .EN(na183_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1048_2_i) );
// C_///AND/D      x112y67     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1049_4 ( .OUT(na1049_2_i), .IN1(na2408_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1049_5 ( .OUT(na1049_2), .CLK(na2414_1), .EN(na183_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1049_2_i) );
// C_///AND/D      x121y81     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1050_4 ( .OUT(na1050_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1050_5 ( .OUT(na1050_2), .CLK(na2414_1), .EN(na183_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1050_2_i) );
// C_AND/D///      x139y72     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1051_1 ( .OUT(na1051_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1051_2 ( .OUT(na1051_1), .CLK(na2414_1), .EN(na183_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1051_1_i) );
// C_///AND/D      x138y31     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1052_4 ( .OUT(na1052_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1052_5 ( .OUT(na1052_2), .CLK(na2414_1), .EN(na184_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1052_2_i) );
// C_AND/D///      x125y38     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1053_1 ( .OUT(na1053_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1053_2 ( .OUT(na1053_1), .CLK(na2414_1), .EN(na184_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1053_1_i) );
// C_///AND/D      x111y45     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1054_4 ( .OUT(na1054_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1054_5 ( .OUT(na1054_2), .CLK(na2414_1), .EN(na184_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1054_2_i) );
// C_AND/D///      x119y49     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1055_1 ( .OUT(na1055_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1055_2 ( .OUT(na1055_1), .CLK(na2414_1), .EN(na184_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1055_1_i) );
// C_AND/D///      x115y51     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1056_1 ( .OUT(na1056_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2405_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1056_2 ( .OUT(na1056_1), .CLK(na2414_1), .EN(na184_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1056_1_i) );
// C_AND/D///      x120y57     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1057_1 ( .OUT(na1057_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1057_2 ( .OUT(na1057_1), .CLK(na2414_1), .EN(na184_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1057_1_i) );
// C_///AND/D      x119y65     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1058_4 ( .OUT(na1058_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1058_5 ( .OUT(na1058_2), .CLK(na2414_1), .EN(na184_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1058_2_i) );
// C_AND/D///      x114y68     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1059_1 ( .OUT(na1059_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1059_2 ( .OUT(na1059_1), .CLK(na2414_1), .EN(na184_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1059_1_i) );
// C_///AND/D      x127y78     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1060_4 ( .OUT(na1060_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1060_5 ( .OUT(na1060_2), .CLK(na2414_1), .EN(na184_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1060_2_i) );
// C_AND/D///      x141y71     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1061_1 ( .OUT(na1061_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1061_2 ( .OUT(na1061_1), .CLK(na2414_1), .EN(na184_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1061_1_i) );
// C_///AND/D      x137y32     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1062_4 ( .OUT(na1062_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1062_5 ( .OUT(na1062_2), .CLK(na2414_1), .EN(na185_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1062_2_i) );
// C_///AND/D      x124y37     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1063_4 ( .OUT(na1063_2_i), .IN1(na2402_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1063_5 ( .OUT(na1063_2), .CLK(na2414_1), .EN(na185_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1063_2_i) );
// C_///AND/D      x116y48     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1064_4 ( .OUT(na1064_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1064_5 ( .OUT(na1064_2), .CLK(na2414_1), .EN(na185_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1064_2_i) );
// C_AND/D///      x120y50     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1065_1 ( .OUT(na1065_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1065_2 ( .OUT(na1065_1), .CLK(na2414_1), .EN(na185_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1065_1_i) );
// C_///AND/D      x120y52     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1066_4 ( .OUT(na1066_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1066_5 ( .OUT(na1066_2), .CLK(na2414_1), .EN(na185_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1066_2_i) );
// C_AND/D///      x119y60     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1067_1 ( .OUT(na1067_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1067_2 ( .OUT(na1067_1), .CLK(na2414_1), .EN(na185_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1067_1_i) );
// C_///AND/D      x122y66     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1068_4 ( .OUT(na1068_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1068_5 ( .OUT(na1068_2), .CLK(na2414_1), .EN(na185_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1068_2_i) );
// C_AND/D///      x115y67     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1069_1 ( .OUT(na1069_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1069_2 ( .OUT(na1069_1), .CLK(na2414_1), .EN(na185_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1069_1_i) );
// C_AND/D///      x116y83     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1070_1 ( .OUT(na1070_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2409_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1070_2 ( .OUT(na1070_1), .CLK(na2414_1), .EN(na185_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1070_1_i) );
// C_AND/D///      x140y72     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1071_1 ( .OUT(na1071_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1071_2 ( .OUT(na1071_1), .CLK(na2414_1), .EN(na185_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1071_1_i) );
// C_///AND/D      x145y30     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1072_4 ( .OUT(na1072_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1072_5 ( .OUT(na1072_2), .CLK(na2414_1), .EN(na180_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1072_2_i) );
// C_AND/D///      x121y38     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1073_1 ( .OUT(na1073_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1073_2 ( .OUT(na1073_1), .CLK(na2414_1), .EN(na180_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1073_1_i) );
// C_///AND/D      x112y43     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1074_4 ( .OUT(na1074_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1074_5 ( .OUT(na1074_2), .CLK(na2414_1), .EN(na180_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1074_2_i) );
// C_AND/D///      x120y48     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1075_1 ( .OUT(na1075_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1075_2 ( .OUT(na1075_1), .CLK(na2414_1), .EN(na180_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1075_1_i) );
// C_///AND/D      x119y58     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1076_4 ( .OUT(na1076_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1076_5 ( .OUT(na1076_2), .CLK(na2414_1), .EN(na180_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1076_2_i) );
// C_///AND/D      x121y60     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1077_4 ( .OUT(na1077_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2406_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1077_5 ( .OUT(na1077_2), .CLK(na2414_1), .EN(na180_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1077_2_i) );
// C_///AND/D      x119y73     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1078_4 ( .OUT(na1078_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1078_5 ( .OUT(na1078_2), .CLK(na2414_1), .EN(na180_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1078_2_i) );
// C_AND/D///      x111y72     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1079_1 ( .OUT(na1079_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1079_2 ( .OUT(na1079_1), .CLK(na2414_1), .EN(na180_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1079_1_i) );
// C_///AND/D      x119y74     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1080_4 ( .OUT(na1080_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1080_5 ( .OUT(na1080_2), .CLK(na2414_1), .EN(na180_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1080_2_i) );
// C_AND/D///      x137y71     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1081_1 ( .OUT(na1081_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1081_2 ( .OUT(na1081_1), .CLK(na2414_1), .EN(na180_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1081_1_i) );
// C_///AND/D      x132y33     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1082_4 ( .OUT(na1082_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1082_5 ( .OUT(na1082_2), .CLK(na2414_1), .EN(na203_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1082_2_i) );
// C_AND/D///      x130y33     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1083_1 ( .OUT(na1083_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1083_2 ( .OUT(na1083_1), .CLK(na2414_1), .EN(na203_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1083_1_i) );
// C_AND/D///      x128y39     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1084_1 ( .OUT(na1084_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2403_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1084_2 ( .OUT(na1084_1), .CLK(na2414_1), .EN(na203_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1084_1_i) );
// C_AND/D///      x138y44     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1085_1 ( .OUT(na1085_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1085_2 ( .OUT(na1085_1), .CLK(na2414_1), .EN(na203_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1085_1_i) );
// C_///AND/D      x129y51     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1086_4 ( .OUT(na1086_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1086_5 ( .OUT(na1086_2), .CLK(na2414_1), .EN(na203_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1086_2_i) );
// C_AND/D///      x121y58     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1087_1 ( .OUT(na1087_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1087_2 ( .OUT(na1087_1), .CLK(na2414_1), .EN(na203_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1087_1_i) );
// C_///AND/D      x121y70     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1088_4 ( .OUT(na1088_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1088_5 ( .OUT(na1088_2), .CLK(na2414_1), .EN(na203_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1088_2_i) );
// C_AND/D///      x117y72     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1089_1 ( .OUT(na1089_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1089_2 ( .OUT(na1089_1), .CLK(na2414_1), .EN(na203_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1089_1_i) );
// C_///AND/D      x136y78     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1090_4 ( .OUT(na1090_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1090_5 ( .OUT(na1090_2), .CLK(na2414_1), .EN(na203_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1090_2_i) );
// C_///AND/D      x133y82     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1091_4 ( .OUT(na1091_2_i), .IN1(1'b1), .IN2(na2410_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1091_5 ( .OUT(na1091_2), .CLK(na2414_1), .EN(na203_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1091_2_i) );
// C_///AND/D      x129y37     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1092_4 ( .OUT(na1092_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1092_5 ( .OUT(na1092_2), .CLK(na2414_1), .EN(na189_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1092_2_i) );
// C_AND/D///      x126y38     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1093_1 ( .OUT(na1093_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1093_2 ( .OUT(na1093_1), .CLK(na2414_1), .EN(na189_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1093_1_i) );
// C_///AND/D      x122y39     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1094_4 ( .OUT(na1094_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1094_5 ( .OUT(na1094_2), .CLK(na2414_1), .EN(na189_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1094_2_i) );
// C_AND/D///      x136y40     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1095_1 ( .OUT(na1095_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1095_2 ( .OUT(na1095_1), .CLK(na2414_1), .EN(na189_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1095_1_i) );
// C_///AND/D      x127y52     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1096_4 ( .OUT(na1096_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1096_5 ( .OUT(na1096_2), .CLK(na2414_1), .EN(na189_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1096_2_i) );
// C_AND/D///      x122y62     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1097_1 ( .OUT(na1097_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1097_2 ( .OUT(na1097_1), .CLK(na2414_1), .EN(na189_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1097_1_i) );
// C_AND/D///      x119y67     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1098_1 ( .OUT(na1098_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2407_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1098_2 ( .OUT(na1098_1), .CLK(na2414_1), .EN(na189_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1098_1_i) );
// C_AND/D///      x115y70     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1099_1 ( .OUT(na1099_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1099_2 ( .OUT(na1099_1), .CLK(na2414_1), .EN(na189_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1099_1_i) );
// C_///AND/D      x127y74     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1100_4 ( .OUT(na1100_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1100_5 ( .OUT(na1100_2), .CLK(na2414_1), .EN(na189_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1100_2_i) );
// C_AND/D///      x127y79     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1101_1 ( .OUT(na1101_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1101_2 ( .OUT(na1101_1), .CLK(na2414_1), .EN(na189_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1101_1_i) );
// C_///AND/D      x132y38     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1102_4 ( .OUT(na1102_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1102_5 ( .OUT(na1102_2), .CLK(na2414_1), .EN(na190_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1102_2_i) );
// C_AND/D///      x127y37     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1103_1 ( .OUT(na1103_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1103_2 ( .OUT(na1103_1), .CLK(na2414_1), .EN(na190_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1103_1_i) );
// C_///AND/D      x123y42     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1104_4 ( .OUT(na1104_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1104_5 ( .OUT(na1104_2), .CLK(na2414_1), .EN(na190_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1104_2_i) );
// C_///AND/D      x133y43     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1105_4 ( .OUT(na1105_2_i), .IN1(1'b1), .IN2(na2404_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1105_5 ( .OUT(na1105_2), .CLK(na2414_1), .EN(na190_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1105_2_i) );
// C_///AND/D      x126y51     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1106_4 ( .OUT(na1106_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1106_5 ( .OUT(na1106_2), .CLK(na2414_1), .EN(na190_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1106_2_i) );
// C_AND/D///      x121y61     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1107_1 ( .OUT(na1107_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1107_2 ( .OUT(na1107_1), .CLK(na2414_1), .EN(na190_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1107_1_i) );
// C_///AND/D      x122y74     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1108_4 ( .OUT(na1108_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1108_5 ( .OUT(na1108_2), .CLK(na2414_1), .EN(na190_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1108_2_i) );
// C_AND/D///      x120y69     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1109_1 ( .OUT(na1109_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1109_2 ( .OUT(na1109_1), .CLK(na2414_1), .EN(na190_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1109_1_i) );
// C_///AND/D      x132y73     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1110_4 ( .OUT(na1110_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1110_5 ( .OUT(na1110_2), .CLK(na2414_1), .EN(na190_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1110_2_i) );
// C_AND/D///      x128y80     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1111_1 ( .OUT(na1111_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1111_2 ( .OUT(na1111_1), .CLK(na2414_1), .EN(na190_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1111_1_i) );
// C_AND/D///      x126y33     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1112_1 ( .OUT(na1112_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2401_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1112_2 ( .OUT(na1112_1), .CLK(na2414_1), .EN(na191_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1112_1_i) );
// C_AND/D///      x129y40     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1113_1 ( .OUT(na1113_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1113_2 ( .OUT(na1113_1), .CLK(na2414_1), .EN(na191_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1113_1_i) );
// C_///AND/D      x121y37     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1114_4 ( .OUT(na1114_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1114_5 ( .OUT(na1114_2), .CLK(na2414_1), .EN(na191_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1114_2_i) );
// C_AND/D///      x135y42     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1115_1 ( .OUT(na1115_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1115_2 ( .OUT(na1115_1), .CLK(na2414_1), .EN(na191_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1115_1_i) );
// C_///AND/D      x126y50     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1116_4 ( .OUT(na1116_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1116_5 ( .OUT(na1116_2), .CLK(na2414_1), .EN(na191_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1116_2_i) );
// C_AND/D///      x121y64     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1117_1 ( .OUT(na1117_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1117_2 ( .OUT(na1117_1), .CLK(na2414_1), .EN(na191_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1117_1_i) );
// C_///AND/D      x124y71     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1118_4 ( .OUT(na1118_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1118_5 ( .OUT(na1118_2), .CLK(na2414_1), .EN(na191_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1118_2_i) );
// C_///AND/D      x124y74     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1119_4 ( .OUT(na1119_2_i), .IN1(na2408_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1119_5 ( .OUT(na1119_2), .CLK(na2414_1), .EN(na191_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1119_2_i) );
// C_///AND/D      x126y76     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1120_4 ( .OUT(na1120_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1120_5 ( .OUT(na1120_2), .CLK(na2414_1), .EN(na191_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1120_2_i) );
// C_AND/D///      x130y79     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1121_1 ( .OUT(na1121_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1121_2 ( .OUT(na1121_1), .CLK(na2414_1), .EN(na191_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1121_1_i) );
// C_///AND/D      x127y34     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1122_4 ( .OUT(na1122_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1122_5 ( .OUT(na1122_2), .CLK(na2414_1), .EN(na192_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1122_2_i) );
// C_AND/D///      x128y38     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1123_1 ( .OUT(na1123_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1123_2 ( .OUT(na1123_1), .CLK(na2414_1), .EN(na192_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1123_1_i) );
// C_///AND/D      x122y36     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1124_4 ( .OUT(na1124_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1124_5 ( .OUT(na1124_2), .CLK(na2414_1), .EN(na192_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1124_2_i) );
// C_AND/D///      x131y43     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1125_1 ( .OUT(na1125_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1125_2 ( .OUT(na1125_1), .CLK(na2414_1), .EN(na192_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1125_1_i) );
// C_AND/D///      x134y57     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1126_1 ( .OUT(na1126_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2405_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1126_2 ( .OUT(na1126_1), .CLK(na2414_1), .EN(na192_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1126_1_i) );
// C_AND/D///      x123y65     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1127_1 ( .OUT(na1127_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1127_2 ( .OUT(na1127_1), .CLK(na2414_1), .EN(na192_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1127_1_i) );
// C_///AND/D      x126y78     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1128_4 ( .OUT(na1128_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1128_5 ( .OUT(na1128_2), .CLK(na2414_1), .EN(na192_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1128_2_i) );
// C_AND/D///      x117y73     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1129_1 ( .OUT(na1129_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1129_2 ( .OUT(na1129_1), .CLK(na2414_1), .EN(na192_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1129_1_i) );
// C_///AND/D      x134y67     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1130_4 ( .OUT(na1130_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1130_5 ( .OUT(na1130_2), .CLK(na2414_1), .EN(na192_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1130_2_i) );
// C_AND/D///      x127y82     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1131_1 ( .OUT(na1131_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1131_2 ( .OUT(na1131_1), .CLK(na2414_1), .EN(na192_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1131_1_i) );
// C_///AND/D      x129y35     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1132_4 ( .OUT(na1132_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1132_5 ( .OUT(na1132_2), .CLK(na2414_1), .EN(na193_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1132_2_i) );
// C_///AND/D      x134y39     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1133_4 ( .OUT(na1133_2_i), .IN1(na2402_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1133_5 ( .OUT(na1133_2), .CLK(na2414_1), .EN(na193_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1133_2_i) );
// C_///AND/D      x124y33     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1134_4 ( .OUT(na1134_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1134_5 ( .OUT(na1134_2), .CLK(na2414_1), .EN(na193_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1134_2_i) );
// C_AND/D///      x133y46     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1135_1 ( .OUT(na1135_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1135_2 ( .OUT(na1135_1), .CLK(na2414_1), .EN(na193_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1135_1_i) );
// C_///AND/D      x126y56     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1136_4 ( .OUT(na1136_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1136_5 ( .OUT(na1136_2), .CLK(na2414_1), .EN(na193_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1136_2_i) );
// C_AND/D///      x125y66     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1137_1 ( .OUT(na1137_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1137_2 ( .OUT(na1137_1), .CLK(na2414_1), .EN(na193_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1137_1_i) );
// C_///AND/D      x122y75     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1138_4 ( .OUT(na1138_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1138_5 ( .OUT(na1138_2), .CLK(na2414_1), .EN(na193_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1138_2_i) );
// C_AND/D///      x115y74     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1139_1 ( .OUT(na1139_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1139_2 ( .OUT(na1139_1), .CLK(na2414_1), .EN(na193_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1139_1_i) );
// C_AND/D///      x128y72     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1140_1 ( .OUT(na1140_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2409_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1140_2 ( .OUT(na1140_1), .CLK(na2414_1), .EN(na193_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1140_1_i) );
// C_AND/D///      x131y81     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1141_1 ( .OUT(na1141_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1141_2 ( .OUT(na1141_1), .CLK(na2414_1), .EN(na193_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1141_1_i) );
// C_///AND/D      x126y34     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1142_4 ( .OUT(na1142_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1142_5 ( .OUT(na1142_2), .CLK(na2414_1), .EN(na194_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1142_2_i) );
// C_AND/D///      x129y38     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1143_1 ( .OUT(na1143_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1143_2 ( .OUT(na1143_1), .CLK(na2414_1), .EN(na194_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1143_1_i) );
// C_///AND/D      x123y36     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1144_4 ( .OUT(na1144_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1144_5 ( .OUT(na1144_2), .CLK(na2414_1), .EN(na194_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1144_2_i) );
// C_AND/D///      x136y45     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1145_1 ( .OUT(na1145_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1145_2 ( .OUT(na1145_1), .CLK(na2414_1), .EN(na194_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1145_1_i) );
// C_///AND/D      x129y55     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1146_4 ( .OUT(na1146_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1146_5 ( .OUT(na1146_2), .CLK(na2414_1), .EN(na194_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1146_2_i) );
// C_///AND/D      x126y65     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1147_4 ( .OUT(na1147_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2406_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1147_5 ( .OUT(na1147_2), .CLK(na2414_1), .EN(na194_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1147_2_i) );
// C_///AND/D      x121y76     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1148_4 ( .OUT(na1148_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1148_5 ( .OUT(na1148_2), .CLK(na2414_1), .EN(na194_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1148_2_i) );
// C_AND/D///      x120y73     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1149_1 ( .OUT(na1149_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1149_2 ( .OUT(na1149_1), .CLK(na2414_1), .EN(na194_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1149_1_i) );
// C_///AND/D      x133y73     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1150_4 ( .OUT(na1150_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1150_5 ( .OUT(na1150_2), .CLK(na2414_1), .EN(na194_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1150_2_i) );
// C_AND/D///      x130y82     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1151_1 ( .OUT(na1151_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1151_2 ( .OUT(na1151_1), .CLK(na2414_1), .EN(na194_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1151_1_i) );
// C_///AND/D      x132y35     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1152_4 ( .OUT(na1152_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1152_5 ( .OUT(na1152_2), .CLK(na2414_1), .EN(na195_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1152_2_i) );
// C_AND/D///      x127y39     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1153_1 ( .OUT(na1153_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1153_2 ( .OUT(na1153_1), .CLK(na2414_1), .EN(na195_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1153_1_i) );
// C_AND/D///      x125y33     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1154_1 ( .OUT(na1154_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2403_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1154_2 ( .OUT(na1154_1), .CLK(na2414_1), .EN(na195_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1154_1_i) );
// C_AND/D///      x134y46     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1155_1 ( .OUT(na1155_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1155_2 ( .OUT(na1155_1), .CLK(na2414_1), .EN(na195_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1155_1_i) );
// C_///AND/D      x127y54     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1156_4 ( .OUT(na1156_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1156_5 ( .OUT(na1156_2), .CLK(na2414_1), .EN(na195_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1156_2_i) );
// C_AND/D///      x128y66     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1157_1 ( .OUT(na1157_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1157_2 ( .OUT(na1157_1), .CLK(na2414_1), .EN(na195_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1157_1_i) );
// C_///AND/D      x121y77     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1158_4 ( .OUT(na1158_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1158_5 ( .OUT(na1158_2), .CLK(na2414_1), .EN(na195_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1158_2_i) );
// C_AND/D///      x118y76     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1159_1 ( .OUT(na1159_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1159_2 ( .OUT(na1159_1), .CLK(na2414_1), .EN(na195_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1159_1_i) );
// C_///AND/D      x131y74     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1160_4 ( .OUT(na1160_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1160_5 ( .OUT(na1160_2), .CLK(na2414_1), .EN(na195_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1160_2_i) );
// C_///AND/D      x130y83     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1161_4 ( .OUT(na1161_2_i), .IN1(1'b1), .IN2(na2410_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1161_5 ( .OUT(na1161_2), .CLK(na2414_1), .EN(na195_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1161_2_i) );
// C_///AND/D      x124y32     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1162_4 ( .OUT(na1162_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1162_5 ( .OUT(na1162_2), .CLK(na2414_1), .EN(na196_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1162_2_i) );
// C_AND/D///      x127y35     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1163_1 ( .OUT(na1163_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1163_2 ( .OUT(na1163_1), .CLK(na2414_1), .EN(na196_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1163_1_i) );
// C_///AND/D      x126y35     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1164_4 ( .OUT(na1164_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1164_5 ( .OUT(na1164_2), .CLK(na2414_1), .EN(na196_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1164_2_i) );
// C_AND/D///      x131y46     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1165_1 ( .OUT(na1165_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1165_2 ( .OUT(na1165_1), .CLK(na2414_1), .EN(na196_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1165_1_i) );
// C_///AND/D      x126y57     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1166_4 ( .OUT(na1166_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1166_5 ( .OUT(na1166_2), .CLK(na2414_1), .EN(na196_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1166_2_i) );
// C_AND/D///      x126y61     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1167_1 ( .OUT(na1167_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1167_2 ( .OUT(na1167_1), .CLK(na2414_1), .EN(na196_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1167_1_i) );
// C_AND/D///      x120y66     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1168_1 ( .OUT(na1168_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2407_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1168_2 ( .OUT(na1168_1), .CLK(na2414_1), .EN(na196_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1168_1_i) );
// C_AND/D///      x120y71     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1169_1 ( .OUT(na1169_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1169_2 ( .OUT(na1169_1), .CLK(na2414_1), .EN(na196_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1169_1_i) );
// C_///AND/D      x129y77     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1170_4 ( .OUT(na1170_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1170_5 ( .OUT(na1170_2), .CLK(na2414_1), .EN(na196_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1170_2_i) );
// C_AND/D///      x127y75     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1171_1 ( .OUT(na1171_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1171_2 ( .OUT(na1171_1), .CLK(na2414_1), .EN(na196_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1171_1_i) );
// C_///AND/D      x127y38     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1172_4 ( .OUT(na1172_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1172_5 ( .OUT(na1172_2), .CLK(na2414_1), .EN(na187_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1172_2_i) );
// C_AND/D///      x130y39     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1173_1 ( .OUT(na1173_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1173_2 ( .OUT(na1173_1), .CLK(na2414_1), .EN(na187_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1173_1_i) );
// C_///AND/D      x128y40     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1174_4 ( .OUT(na1174_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1174_5 ( .OUT(na1174_2), .CLK(na2414_1), .EN(na187_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1174_2_i) );
// C_///AND/D      x138y43     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1175_4 ( .OUT(na1175_2_i), .IN1(1'b1), .IN2(na2404_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1175_5 ( .OUT(na1175_2), .CLK(na2414_1), .EN(na187_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1175_2_i) );
// C_///AND/D      x133y47     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1176_4 ( .OUT(na1176_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1176_5 ( .OUT(na1176_2), .CLK(na2414_1), .EN(na187_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1176_2_i) );
// C_AND/D///      x122y63     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1177_1 ( .OUT(na1177_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1177_2 ( .OUT(na1177_1), .CLK(na2414_1), .EN(na187_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1177_1_i) );
// C_///AND/D      x121y72     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1178_4 ( .OUT(na1178_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1178_5 ( .OUT(na1178_2), .CLK(na2414_1), .EN(na187_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1178_2_i) );
// C_AND/D///      x115y71     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1179_1 ( .OUT(na1179_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1179_2 ( .OUT(na1179_1), .CLK(na2414_1), .EN(na187_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1179_1_i) );
// C_///AND/D      x129y75     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1180_4 ( .OUT(na1180_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1180_5 ( .OUT(na1180_2), .CLK(na2414_1), .EN(na187_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1180_2_i) );
// C_AND/D///      x129y80     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1181_1 ( .OUT(na1181_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1181_2 ( .OUT(na1181_1), .CLK(na2414_1), .EN(na187_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1181_1_i) );
// C_AND/D///      x129y32     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1182_1 ( .OUT(na1182_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2401_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1182_2 ( .OUT(na1182_1), .CLK(na2414_1), .EN(na198_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1182_1_i) );
// C_AND/D///      x130y35     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1183_1 ( .OUT(na1183_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1183_2 ( .OUT(na1183_1), .CLK(na2414_1), .EN(na198_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1183_1_i) );
// C_///AND/D      x129y39     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1184_4 ( .OUT(na1184_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1184_5 ( .OUT(na1184_2), .CLK(na2414_1), .EN(na198_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1184_2_i) );
// C_AND/D///      x130y46     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1185_1 ( .OUT(na1185_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1185_2 ( .OUT(na1185_1), .CLK(na2414_1), .EN(na198_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1185_1_i) );
// C_///AND/D      x129y57     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1186_4 ( .OUT(na1186_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1186_5 ( .OUT(na1186_2), .CLK(na2414_1), .EN(na198_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1186_2_i) );
// C_AND/D///      x123y61     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1187_1 ( .OUT(na1187_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1187_2 ( .OUT(na1187_1), .CLK(na2414_1), .EN(na198_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1187_1_i) );
// C_///AND/D      x123y70     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1188_4 ( .OUT(na1188_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1188_5 ( .OUT(na1188_2), .CLK(na2414_1), .EN(na198_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1188_2_i) );
// C_///AND/D      x117y71     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1189_4 ( .OUT(na1189_2_i), .IN1(na2408_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1189_5 ( .OUT(na1189_2), .CLK(na2414_1), .EN(na198_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1189_2_i) );
// C_///AND/D      x132y79     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1190_4 ( .OUT(na1190_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1190_5 ( .OUT(na1190_2), .CLK(na2414_1), .EN(na198_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1190_2_i) );
// C_AND/D///      x128y77     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1191_1 ( .OUT(na1191_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1191_2 ( .OUT(na1191_1), .CLK(na2414_1), .EN(na198_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1191_1_i) );
// C_///AND/D      x131y33     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1192_4 ( .OUT(na1192_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1192_5 ( .OUT(na1192_2), .CLK(na2414_1), .EN(na199_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1192_2_i) );
// C_AND/D///      x128y34     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1193_1 ( .OUT(na1193_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1193_2 ( .OUT(na1193_1), .CLK(na2414_1), .EN(na199_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1193_1_i) );
// C_///AND/D      x127y40     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1194_4 ( .OUT(na1194_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1194_5 ( .OUT(na1194_2), .CLK(na2414_1), .EN(na199_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1194_2_i) );
// C_AND/D///      x132y45     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1195_1 ( .OUT(na1195_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1195_2 ( .OUT(na1195_1), .CLK(na2414_1), .EN(na199_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1195_1_i) );
// C_AND/D///      x131y58     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1196_1 ( .OUT(na1196_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2405_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1196_2 ( .OUT(na1196_1), .CLK(na2414_1), .EN(na199_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1196_1_i) );
// C_AND/D///      x125y62     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1197_1 ( .OUT(na1197_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1197_2 ( .OUT(na1197_1), .CLK(na2414_1), .EN(na199_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1197_1_i) );
// C_///AND/D      x125y69     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1198_4 ( .OUT(na1198_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1198_5 ( .OUT(na1198_2), .CLK(na2414_1), .EN(na199_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1198_2_i) );
// C_AND/D///      x119y72     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1199_1 ( .OUT(na1199_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1199_2 ( .OUT(na1199_1), .CLK(na2414_1), .EN(na199_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1199_1_i) );
// C_///AND/D      x132y82     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1200_4 ( .OUT(na1200_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1200_5 ( .OUT(na1200_2), .CLK(na2414_1), .EN(na199_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1200_2_i) );
// C_AND/D///      x130y78     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1201_1 ( .OUT(na1201_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1201_2 ( .OUT(na1201_1), .CLK(na2414_1), .EN(na199_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1201_1_i) );
// C_///AND/D      x131y36     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1202_4 ( .OUT(na1202_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1202_5 ( .OUT(na1202_2), .CLK(na2414_1), .EN(na200_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1202_2_i) );
// C_///AND/D      x131y38     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1203_4 ( .OUT(na1203_2_i), .IN1(na2402_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1203_5 ( .OUT(na1203_2), .CLK(na2414_1), .EN(na200_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1203_2_i) );
// C_///AND/D      x127y42     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1204_4 ( .OUT(na1204_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1204_5 ( .OUT(na1204_2), .CLK(na2414_1), .EN(na200_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1204_2_i) );
// C_AND/D///      x135y45     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1205_1 ( .OUT(na1205_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1205_2 ( .OUT(na1205_1), .CLK(na2414_1), .EN(na200_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1205_1_i) );
// C_///AND/D      x132y52     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1206_4 ( .OUT(na1206_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1206_5 ( .OUT(na1206_2), .CLK(na2414_1), .EN(na200_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1206_2_i) );
// C_AND/D///      x122y57     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1207_1 ( .OUT(na1207_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1207_2 ( .OUT(na1207_1), .CLK(na2414_1), .EN(na200_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1207_1_i) );
// C_///AND/D      x124y73     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1208_4 ( .OUT(na1208_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1208_5 ( .OUT(na1208_2), .CLK(na2414_1), .EN(na200_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1208_2_i) );
// C_AND/D///      x118y71     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1209_1 ( .OUT(na1209_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1209_2 ( .OUT(na1209_1), .CLK(na2414_1), .EN(na200_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1209_1_i) );
// C_AND/D///      x129y73     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1210_1 ( .OUT(na1210_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2409_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1210_2 ( .OUT(na1210_1), .CLK(na2414_1), .EN(na200_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1210_1_i) );
// C_AND/D///      x126y81     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1211_1 ( .OUT(na1211_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1211_2 ( .OUT(na1211_1), .CLK(na2414_1), .EN(na200_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1211_1_i) );
// C_///AND/D      x133y37     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1212_4 ( .OUT(na1212_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1212_5 ( .OUT(na1212_2), .CLK(na2414_1), .EN(na201_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1212_2_i) );
// C_AND/D///      x129y33     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1213_1 ( .OUT(na1213_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1213_2 ( .OUT(na1213_1), .CLK(na2414_1), .EN(na201_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1213_1_i) );
// C_///AND/D      x131y39     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1214_4 ( .OUT(na1214_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1214_5 ( .OUT(na1214_2), .CLK(na2414_1), .EN(na201_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1214_2_i) );
// C_AND/D///      x135y46     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1215_1 ( .OUT(na1215_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1215_2 ( .OUT(na1215_1), .CLK(na2414_1), .EN(na201_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1215_1_i) );
// C_///AND/D      x132y53     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1216_4 ( .OUT(na1216_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1216_5 ( .OUT(na1216_2), .CLK(na2414_1), .EN(na201_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1216_2_i) );
// C_///AND/D      x124y64     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1217_4 ( .OUT(na1217_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2406_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1217_5 ( .OUT(na1217_2), .CLK(na2414_1), .EN(na201_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1217_2_i) );
// C_///AND/D      x126y72     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1218_4 ( .OUT(na1218_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1218_5 ( .OUT(na1218_2), .CLK(na2414_1), .EN(na201_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1218_2_i) );
// C_AND/D///      x116y74     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1219_1 ( .OUT(na1219_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1219_2 ( .OUT(na1219_1), .CLK(na2414_1), .EN(na201_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1219_1_i) );
// C_///AND/D      x131y80     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1220_4 ( .OUT(na1220_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1220_5 ( .OUT(na1220_2), .CLK(na2414_1), .EN(na201_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1220_2_i) );
// C_AND/D///      x126y82     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1221_1 ( .OUT(na1221_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1221_2 ( .OUT(na1221_1), .CLK(na2414_1), .EN(na201_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1221_1_i) );
// C_///AND/D      x132y30     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1222_4 ( .OUT(na1222_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1222_5 ( .OUT(na1222_2), .CLK(na2414_1), .EN(na202_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1222_2_i) );
// C_AND/D///      x130y34     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1223_1 ( .OUT(na1223_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1223_2 ( .OUT(na1223_1), .CLK(na2414_1), .EN(na202_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1223_1_i) );
// C_AND/D///      x126y42     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1224_1 ( .OUT(na1224_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2403_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1224_2 ( .OUT(na1224_1), .CLK(na2414_1), .EN(na202_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1224_1_i) );
// C_AND/D///      x138y45     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1225_1 ( .OUT(na1225_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1225_2 ( .OUT(na1225_1), .CLK(na2414_1), .EN(na202_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1225_1_i) );
// C_///AND/D      x133y50     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1226_4 ( .OUT(na1226_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1226_5 ( .OUT(na1226_2), .CLK(na2414_1), .EN(na202_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1226_2_i) );
// C_AND/D///      x121y59     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1227_1 ( .OUT(na1227_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1227_2 ( .OUT(na1227_1), .CLK(na2414_1), .EN(na202_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1227_1_i) );
// C_///AND/D      x121y69     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1228_4 ( .OUT(na1228_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1228_5 ( .OUT(na1228_2), .CLK(na2414_1), .EN(na202_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1228_2_i) );
// C_AND/D///      x115y73     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1229_1 ( .OUT(na1229_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1229_2 ( .OUT(na1229_1), .CLK(na2414_1), .EN(na202_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1229_1_i) );
// C_///AND/D      x132y77     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1230_4 ( .OUT(na1230_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1230_5 ( .OUT(na1230_2), .CLK(na2414_1), .EN(na202_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1230_2_i) );
// C_///AND/D      x129y83     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1231_4 ( .OUT(na1231_2_i), .IN1(1'b1), .IN2(na2410_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1231_5 ( .OUT(na1231_2), .CLK(na2414_1), .EN(na202_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1231_2_i) );
// C_///AND/D      x128y33     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1232_4 ( .OUT(na1232_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1232_5 ( .OUT(na1232_2), .CLK(na2414_1), .EN(na197_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1232_2_i) );
// C_AND/D///      x129y36     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1233_1 ( .OUT(na1233_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1233_2 ( .OUT(na1233_1), .CLK(na2414_1), .EN(na197_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1233_1_i) );
// C_///AND/D      x132y40     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1234_4 ( .OUT(na1234_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1234_5 ( .OUT(na1234_2), .CLK(na2414_1), .EN(na197_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1234_2_i) );
// C_AND/D///      x131y47     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1235_1 ( .OUT(na1235_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1235_2 ( .OUT(na1235_1), .CLK(na2414_1), .EN(na197_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1235_1_i) );
// C_///AND/D      x132y56     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1236_4 ( .OUT(na1236_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1236_5 ( .OUT(na1236_2), .CLK(na2414_1), .EN(na197_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1236_2_i) );
// C_AND/D///      x128y64     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1237_1 ( .OUT(na1237_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1237_2 ( .OUT(na1237_1), .CLK(na2414_1), .EN(na197_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1237_1_i) );
// C_AND/D///      x120y67     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1238_1 ( .OUT(na1238_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2407_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1238_2 ( .OUT(na1238_1), .CLK(na2414_1), .EN(na197_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1238_1_i) );
// C_AND/D///      x120y72     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1239_1 ( .OUT(na1239_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1239_2 ( .OUT(na1239_1), .CLK(na2414_1), .EN(na197_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1239_1_i) );
// C_///AND/D      x129y78     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1240_4 ( .OUT(na1240_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1240_5 ( .OUT(na1240_2), .CLK(na2414_1), .EN(na197_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1240_2_i) );
// C_AND/D///      x129y78     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1241_1 ( .OUT(na1241_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1241_2 ( .OUT(na1241_1), .CLK(na2414_1), .EN(na197_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1241_1_i) );
// C_///AND/D      x147y42     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1242_4 ( .OUT(na1242_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1242_5 ( .OUT(na1242_2), .CLK(na2414_1), .EN(na220_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1242_2_i) );
// C_AND/D///      x131y35     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1243_1 ( .OUT(na1243_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1243_2 ( .OUT(na1243_1), .CLK(na2414_1), .EN(na220_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1243_1_i) );
// C_///AND/D      x145y56     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1244_4 ( .OUT(na1244_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1244_5 ( .OUT(na1244_2), .CLK(na2414_1), .EN(na220_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1244_2_i) );
// C_///AND/D      x136y51     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1245_4 ( .OUT(na1245_2_i), .IN1(1'b1), .IN2(na2404_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1245_5 ( .OUT(na1245_2), .CLK(na2414_1), .EN(na220_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1245_2_i) );
// C_///AND/D      x148y56     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1246_4 ( .OUT(na1246_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1246_5 ( .OUT(na1246_2), .CLK(na2414_1), .EN(na220_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1246_2_i) );
// C_AND/D///      x154y54     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1247_1 ( .OUT(na1247_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1247_2 ( .OUT(na1247_1), .CLK(na2414_1), .EN(na220_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1247_1_i) );
// C_///AND/D      x143y74     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1248_4 ( .OUT(na1248_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1248_5 ( .OUT(na1248_2), .CLK(na2414_1), .EN(na220_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1248_2_i) );
// C_AND/D///      x148y71     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1249_1 ( .OUT(na1249_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1249_2 ( .OUT(na1249_1), .CLK(na2414_1), .EN(na220_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1249_1_i) );
// C_///AND/D      x156y75     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1250_4 ( .OUT(na1250_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1250_5 ( .OUT(na1250_2), .CLK(na2414_1), .EN(na220_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1250_2_i) );
// C_AND/D///      x143y79     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1251_1 ( .OUT(na1251_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1251_2 ( .OUT(na1251_1), .CLK(na2414_1), .EN(na220_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1251_1_i) );
// C_AND/D///      x151y37     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1252_1 ( .OUT(na1252_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2401_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1252_2 ( .OUT(na1252_1), .CLK(na2414_1), .EN(na206_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1252_1_i) );
// C_AND/D///      x130y43     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1253_1 ( .OUT(na1253_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1253_2 ( .OUT(na1253_1), .CLK(na2414_1), .EN(na206_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1253_1_i) );
// C_///AND/D      x148y54     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1254_4 ( .OUT(na1254_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1254_5 ( .OUT(na1254_2), .CLK(na2414_1), .EN(na206_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1254_2_i) );
// C_AND/D///      x134y50     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1255_1 ( .OUT(na1255_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1255_2 ( .OUT(na1255_1), .CLK(na2414_1), .EN(na206_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1255_1_i) );
// C_///AND/D      x149y61     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1256_4 ( .OUT(na1256_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1256_5 ( .OUT(na1256_2), .CLK(na2414_1), .EN(na206_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1256_2_i) );
// C_AND/D///      x152y57     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1257_1 ( .OUT(na1257_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1257_2 ( .OUT(na1257_1), .CLK(na2414_1), .EN(na206_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1257_1_i) );
// C_///AND/D      x144y70     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1258_4 ( .OUT(na1258_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1258_5 ( .OUT(na1258_2), .CLK(na2414_1), .EN(na206_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1258_2_i) );
// C_///AND/D      x151y66     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1259_4 ( .OUT(na1259_2_i), .IN1(na2408_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1259_5 ( .OUT(na1259_2), .CLK(na2414_1), .EN(na206_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1259_2_i) );
// C_///AND/D      x151y70     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1260_4 ( .OUT(na1260_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1260_5 ( .OUT(na1260_2), .CLK(na2414_1), .EN(na206_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1260_2_i) );
// C_AND/D///      x146y77     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1261_1 ( .OUT(na1261_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1261_2 ( .OUT(na1261_1), .CLK(na2414_1), .EN(na206_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1261_1_i) );
// C_///AND/D      x142y44     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1262_4 ( .OUT(na1262_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1262_5 ( .OUT(na1262_2), .CLK(na2414_1), .EN(na207_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1262_2_i) );
// C_AND/D///      x129y44     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1263_1 ( .OUT(na1263_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1263_2 ( .OUT(na1263_1), .CLK(na2414_1), .EN(na207_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1263_1_i) );
// C_///AND/D      x147y55     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1264_4 ( .OUT(na1264_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1264_5 ( .OUT(na1264_2), .CLK(na2414_1), .EN(na207_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1264_2_i) );
// C_AND/D///      x135y49     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1265_1 ( .OUT(na1265_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1265_2 ( .OUT(na1265_1), .CLK(na2414_1), .EN(na207_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1265_1_i) );
// C_AND/D///      x152y50     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1266_1 ( .OUT(na1266_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2405_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1266_2 ( .OUT(na1266_1), .CLK(na2414_1), .EN(na207_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1266_1_i) );
// C_AND/D///      x155y58     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1267_1 ( .OUT(na1267_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1267_2 ( .OUT(na1267_1), .CLK(na2414_1), .EN(na207_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1267_1_i) );
// C_///AND/D      x143y73     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1268_4 ( .OUT(na1268_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1268_5 ( .OUT(na1268_2), .CLK(na2414_1), .EN(na207_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1268_2_i) );
// C_AND/D///      x156y73     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1269_1 ( .OUT(na1269_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1269_2 ( .OUT(na1269_1), .CLK(na2414_1), .EN(na207_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1269_1_i) );
// C_///AND/D      x152y71     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1270_4 ( .OUT(na1270_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1270_5 ( .OUT(na1270_2), .CLK(na2414_1), .EN(na207_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1270_2_i) );
// C_AND/D///      x147y78     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1271_1 ( .OUT(na1271_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1271_2 ( .OUT(na1271_1), .CLK(na2414_1), .EN(na207_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1271_1_i) );
// C_///AND/D      x144y45     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1272_4 ( .OUT(na1272_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1272_5 ( .OUT(na1272_2), .CLK(na2414_1), .EN(na208_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1272_2_i) );
// C_///AND/D      x133y41     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1273_4 ( .OUT(na1273_2_i), .IN1(na2402_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1273_5 ( .OUT(na1273_2), .CLK(na2414_1), .EN(na208_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1273_2_i) );
// C_///AND/D      x151y52     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1274_4 ( .OUT(na1274_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1274_5 ( .OUT(na1274_2), .CLK(na2414_1), .EN(na208_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1274_2_i) );
// C_AND/D///      x137y50     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1275_1 ( .OUT(na1275_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1275_2 ( .OUT(na1275_1), .CLK(na2414_1), .EN(na208_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1275_1_i) );
// C_///AND/D      x152y61     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1276_4 ( .OUT(na1276_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1276_5 ( .OUT(na1276_2), .CLK(na2414_1), .EN(na208_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1276_2_i) );
// C_AND/D///      x153y59     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1277_1 ( .OUT(na1277_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1277_2 ( .OUT(na1277_1), .CLK(na2414_1), .EN(na208_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1277_1_i) );
// C_///AND/D      x141y72     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1278_4 ( .OUT(na1278_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1278_5 ( .OUT(na1278_2), .CLK(na2414_1), .EN(na208_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1278_2_i) );
// C_AND/D///      x154y74     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1279_1 ( .OUT(na1279_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1279_2 ( .OUT(na1279_1), .CLK(na2414_1), .EN(na208_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1279_1_i) );
// C_AND/D///      x154y78     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1280_1 ( .OUT(na1280_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2409_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1280_2 ( .OUT(na1280_1), .CLK(na2414_1), .EN(na208_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1280_1_i) );
// C_AND/D///      x145y79     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1281_1 ( .OUT(na1281_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1281_2 ( .OUT(na1281_1), .CLK(na2414_1), .EN(na208_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1281_1_i) );
// C_///AND/D      x149y40     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1282_4 ( .OUT(na1282_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1282_5 ( .OUT(na1282_2), .CLK(na2414_1), .EN(na209_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1282_2_i) );
// C_AND/D///      x134y38     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1283_1 ( .OUT(na1283_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1283_2 ( .OUT(na1283_1), .CLK(na2414_1), .EN(na209_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1283_1_i) );
// C_///AND/D      x146y55     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1284_4 ( .OUT(na1284_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1284_5 ( .OUT(na1284_2), .CLK(na2414_1), .EN(na209_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1284_2_i) );
// C_AND/D///      x135y50     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1285_1 ( .OUT(na1285_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1285_2 ( .OUT(na1285_1), .CLK(na2414_1), .EN(na209_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1285_1_i) );
// C_///AND/D      x154y65     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1286_4 ( .OUT(na1286_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1286_5 ( .OUT(na1286_2), .CLK(na2414_1), .EN(na209_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1286_2_i) );
// C_///AND/D      x149y63     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1287_4 ( .OUT(na1287_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2406_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1287_5 ( .OUT(na1287_2), .CLK(na2414_1), .EN(na209_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1287_2_i) );
// C_///AND/D      x145y66     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1288_4 ( .OUT(na1288_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1288_5 ( .OUT(na1288_2), .CLK(na2414_1), .EN(na209_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1288_2_i) );
// C_AND/D///      x150y73     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1289_1 ( .OUT(na1289_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1289_2 ( .OUT(na1289_1), .CLK(na2414_1), .EN(na209_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1289_1_i) );
// C_///AND/D      x144y84     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1290_4 ( .OUT(na1290_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1290_5 ( .OUT(na1290_2), .CLK(na2414_1), .EN(na209_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1290_2_i) );
// C_AND/D///      x143y81     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1291_1 ( .OUT(na1291_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1291_2 ( .OUT(na1291_1), .CLK(na2414_1), .EN(na209_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1291_1_i) );
// C_///AND/D      x149y43     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1292_4 ( .OUT(na1292_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1292_5 ( .OUT(na1292_2), .CLK(na2414_1), .EN(na210_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1292_2_i) );
// C_AND/D///      x132y39     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1293_1 ( .OUT(na1293_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1293_2 ( .OUT(na1293_1), .CLK(na2414_1), .EN(na210_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1293_1_i) );
// C_AND/D///      x150y48     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1294_1 ( .OUT(na1294_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2403_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1294_2 ( .OUT(na1294_1), .CLK(na2414_1), .EN(na210_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1294_1_i) );
// C_AND/D///      x137y49     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1295_1 ( .OUT(na1295_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1295_2 ( .OUT(na1295_1), .CLK(na2414_1), .EN(na210_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1295_1_i) );
// C_///AND/D      x156y62     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1296_4 ( .OUT(na1296_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1296_5 ( .OUT(na1296_2), .CLK(na2414_1), .EN(na210_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1296_2_i) );
// C_AND/D///      x151y58     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1297_1 ( .OUT(na1297_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1297_2 ( .OUT(na1297_1), .CLK(na2414_1), .EN(na210_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1297_1_i) );
// C_///AND/D      x147y69     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1298_4 ( .OUT(na1298_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1298_5 ( .OUT(na1298_2), .CLK(na2414_1), .EN(na210_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1298_2_i) );
// C_AND/D///      x150y76     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1299_1 ( .OUT(na1299_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1299_2 ( .OUT(na1299_1), .CLK(na2414_1), .EN(na210_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1299_1_i) );
// C_///AND/D      x146y81     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1300_4 ( .OUT(na1300_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1300_5 ( .OUT(na1300_2), .CLK(na2414_1), .EN(na210_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1300_2_i) );
// C_///AND/D      x141y80     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1301_4 ( .OUT(na1301_2_i), .IN1(1'b1), .IN2(na2410_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1301_5 ( .OUT(na1301_2), .CLK(na2414_1), .EN(na210_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1301_2_i) );
// C_///AND/D      x154y42     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1302_4 ( .OUT(na1302_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1302_5 ( .OUT(na1302_2), .CLK(na2414_1), .EN(na211_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1302_2_i) );
// C_AND/D///      x131y40     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1303_1 ( .OUT(na1303_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1303_2 ( .OUT(na1303_1), .CLK(na2414_1), .EN(na211_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1303_1_i) );
// C_///AND/D      x145y55     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1304_4 ( .OUT(na1304_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1304_5 ( .OUT(na1304_2), .CLK(na2414_1), .EN(na211_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1304_2_i) );
// C_AND/D///      x136y52     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1305_1 ( .OUT(na1305_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1305_2 ( .OUT(na1305_1), .CLK(na2414_1), .EN(na211_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1305_1_i) );
// C_///AND/D      x155y61     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1306_4 ( .OUT(na1306_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1306_5 ( .OUT(na1306_2), .CLK(na2414_1), .EN(na211_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1306_2_i) );
// C_AND/D///      x154y59     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1307_1 ( .OUT(na1307_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1307_2 ( .OUT(na1307_1), .CLK(na2414_1), .EN(na211_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1307_1_i) );
// C_AND/D///      x148y66     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1308_1 ( .OUT(na1308_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2407_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1308_2 ( .OUT(na1308_1), .CLK(na2414_1), .EN(na211_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1308_1_i) );
// C_AND/D///      x147y75     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1309_1 ( .OUT(na1309_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1309_2 ( .OUT(na1309_1), .CLK(na2414_1), .EN(na211_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1309_1_i) );
// C_///AND/D      x147y82     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1310_4 ( .OUT(na1310_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1310_5 ( .OUT(na1310_2), .CLK(na2414_1), .EN(na211_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1310_2_i) );
// C_AND/D///      x140y79     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1311_1 ( .OUT(na1311_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1311_2 ( .OUT(na1311_1), .CLK(na2414_1), .EN(na211_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1311_1_i) );
// C_///AND/D      x152y45     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1312_4 ( .OUT(na1312_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1312_5 ( .OUT(na1312_2), .CLK(na2414_1), .EN(na212_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1312_2_i) );
// C_AND/D///      x135y37     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1313_1 ( .OUT(na1313_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1313_2 ( .OUT(na1313_1), .CLK(na2414_1), .EN(na212_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1313_1_i) );
// C_///AND/D      x147y56     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1314_4 ( .OUT(na1314_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1314_5 ( .OUT(na1314_2), .CLK(na2414_1), .EN(na212_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1314_2_i) );
// C_///AND/D      x132y49     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1315_4 ( .OUT(na1315_2_i), .IN1(1'b1), .IN2(na2404_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1315_5 ( .OUT(na1315_2), .CLK(na2414_1), .EN(na212_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1315_2_i) );
// C_///AND/D      x155y64     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1316_4 ( .OUT(na1316_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1316_5 ( .OUT(na1316_2), .CLK(na2414_1), .EN(na212_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1316_2_i) );
// C_AND/D///      x152y60     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1317_1 ( .OUT(na1317_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1317_2 ( .OUT(na1317_1), .CLK(na2414_1), .EN(na212_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1317_1_i) );
// C_///AND/D      x144y71     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1318_4 ( .OUT(na1318_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1318_5 ( .OUT(na1318_2), .CLK(na2414_1), .EN(na212_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1318_2_i) );
// C_AND/D///      x149y76     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1319_1 ( .OUT(na1319_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1319_2 ( .OUT(na1319_1), .CLK(na2414_1), .EN(na212_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1319_1_i) );
// C_///AND/D      x149y81     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1320_4 ( .OUT(na1320_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1320_5 ( .OUT(na1320_2), .CLK(na2414_1), .EN(na212_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1320_2_i) );
// C_AND/D///      x142y80     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1321_1 ( .OUT(na1321_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1321_2 ( .OUT(na1321_1), .CLK(na2414_1), .EN(na212_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1321_1_i) );
// C_AND/D///      x150y39     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1322_1 ( .OUT(na1322_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2401_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1322_2 ( .OUT(na1322_1), .CLK(na2414_1), .EN(na213_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1322_1_i) );
// C_AND/D///      x134y40     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1323_1 ( .OUT(na1323_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1323_2 ( .OUT(na1323_1), .CLK(na2414_1), .EN(na213_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1323_1_i) );
// C_///AND/D      x141y49     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1324_4 ( .OUT(na1324_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1324_5 ( .OUT(na1324_2), .CLK(na2414_1), .EN(na213_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1324_2_i) );
// C_AND/D///      x137y53     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1325_1 ( .OUT(na1325_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1325_2 ( .OUT(na1325_1), .CLK(na2414_1), .EN(na213_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1325_1_i) );
// C_///AND/D      x150y55     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1326_4 ( .OUT(na1326_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1326_5 ( .OUT(na1326_2), .CLK(na2414_1), .EN(na213_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1326_2_i) );
// C_AND/D///      x156y59     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1327_1 ( .OUT(na1327_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1327_2 ( .OUT(na1327_1), .CLK(na2414_1), .EN(na213_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1327_1_i) );
// C_///AND/D      x147y74     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1328_4 ( .OUT(na1328_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1328_5 ( .OUT(na1328_2), .CLK(na2414_1), .EN(na213_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1328_2_i) );
// C_///AND/D      x153y73     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1329_4 ( .OUT(na1329_2_i), .IN1(na2408_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1329_5 ( .OUT(na1329_2), .CLK(na2414_1), .EN(na213_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1329_2_i) );
// C_///AND/D      x155y67     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1330_4 ( .OUT(na1330_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1330_5 ( .OUT(na1330_2), .CLK(na2414_1), .EN(na213_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1330_2_i) );
// C_AND/D///      x142y75     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1331_1 ( .OUT(na1331_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1331_2 ( .OUT(na1331_1), .CLK(na2414_1), .EN(na213_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1331_1_i) );
// C_///AND/D      x143y50     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1332_4 ( .OUT(na1332_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1332_5 ( .OUT(na1332_2), .CLK(na2414_1), .EN(na204_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1332_2_i) );
// C_AND/D///      x130y44     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1333_1 ( .OUT(na1333_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1333_2 ( .OUT(na1333_1), .CLK(na2414_1), .EN(na204_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1333_1_i) );
// C_///AND/D      x152y51     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1334_4 ( .OUT(na1334_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1334_5 ( .OUT(na1334_2), .CLK(na2414_1), .EN(na204_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1334_2_i) );
// C_AND/D///      x136y53     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1335_1 ( .OUT(na1335_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1335_2 ( .OUT(na1335_1), .CLK(na2414_1), .EN(na204_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1335_1_i) );
// C_AND/D///      x149y52     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1336_1 ( .OUT(na1336_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2405_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1336_2 ( .OUT(na1336_1), .CLK(na2414_1), .EN(na204_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1336_1_i) );
// C_AND/D///      x154y60     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1337_1 ( .OUT(na1337_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1337_2 ( .OUT(na1337_1), .CLK(na2414_1), .EN(na204_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1337_1_i) );
// C_///AND/D      x144y73     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1338_4 ( .OUT(na1338_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1338_5 ( .OUT(na1338_2), .CLK(na2414_1), .EN(na204_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1338_2_i) );
// C_AND/D///      x153y75     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1339_1 ( .OUT(na1339_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1339_2 ( .OUT(na1339_1), .CLK(na2414_1), .EN(na204_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1339_1_i) );
// C_///AND/D      x155y71     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1340_4 ( .OUT(na1340_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1340_5 ( .OUT(na1340_2), .CLK(na2414_1), .EN(na204_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1340_2_i) );
// C_AND/D///      x148y80     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1341_1 ( .OUT(na1341_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1341_2 ( .OUT(na1341_1), .CLK(na2414_1), .EN(na204_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1341_1_i) );
// C_///AND/D      x143y47     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1342_4 ( .OUT(na1342_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1342_5 ( .OUT(na1342_2), .CLK(na2414_1), .EN(na215_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1342_2_i) );
// C_///AND/D      x131y42     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1343_4 ( .OUT(na1343_2_i), .IN1(na2402_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1343_5 ( .OUT(na1343_2), .CLK(na2414_1), .EN(na215_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1343_2_i) );
// C_///AND/D      x146y49     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1344_4 ( .OUT(na1344_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1344_5 ( .OUT(na1344_2), .CLK(na2414_1), .EN(na215_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1344_2_i) );
// C_AND/D///      x136y55     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1345_1 ( .OUT(na1345_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1345_2 ( .OUT(na1345_1), .CLK(na2414_1), .EN(na215_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1345_1_i) );
// C_///AND/D      x149y59     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1346_4 ( .OUT(na1346_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1346_5 ( .OUT(na1346_2), .CLK(na2414_1), .EN(na215_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1346_2_i) );
// C_AND/D///      x153y61     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1347_1 ( .OUT(na1347_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1347_2 ( .OUT(na1347_1), .CLK(na2414_1), .EN(na215_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1347_1_i) );
// C_///AND/D      x148y72     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1348_4 ( .OUT(na1348_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1348_5 ( .OUT(na1348_2), .CLK(na2414_1), .EN(na215_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1348_2_i) );
// C_AND/D///      x150y69     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1349_1 ( .OUT(na1349_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1349_2 ( .OUT(na1349_1), .CLK(na2414_1), .EN(na215_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1349_1_i) );
// C_AND/D///      x154y75     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1350_1 ( .OUT(na1350_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2409_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1350_2 ( .OUT(na1350_1), .CLK(na2414_1), .EN(na215_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1350_1_i) );
// C_AND/D///      x143y77     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1351_1 ( .OUT(na1351_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1351_2 ( .OUT(na1351_1), .CLK(na2414_1), .EN(na215_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1351_1_i) );
// C_///AND/D      x143y46     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1352_4 ( .OUT(na1352_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1352_5 ( .OUT(na1352_2), .CLK(na2414_1), .EN(na216_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1352_2_i) );
// C_AND/D///      x131y41     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1353_1 ( .OUT(na1353_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1353_2 ( .OUT(na1353_1), .CLK(na2414_1), .EN(na216_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1353_1_i) );
// C_///AND/D      x142y46     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1354_4 ( .OUT(na1354_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1354_5 ( .OUT(na1354_2), .CLK(na2414_1), .EN(na216_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1354_2_i) );
// C_AND/D///      x136y56     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1355_1 ( .OUT(na1355_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1355_2 ( .OUT(na1355_1), .CLK(na2414_1), .EN(na216_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1355_1_i) );
// C_///AND/D      x149y58     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1356_4 ( .OUT(na1356_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1356_5 ( .OUT(na1356_2), .CLK(na2414_1), .EN(na216_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1356_2_i) );
// C_///AND/D      x157y64     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1357_4 ( .OUT(na1357_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2406_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1357_5 ( .OUT(na1357_2), .CLK(na2414_1), .EN(na216_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1357_2_i) );
// C_///AND/D      x148y75     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1358_4 ( .OUT(na1358_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1358_5 ( .OUT(na1358_2), .CLK(na2414_1), .EN(na216_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1358_2_i) );
// C_AND/D///      x150y70     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1359_1 ( .OUT(na1359_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1359_2 ( .OUT(na1359_1), .CLK(na2414_1), .EN(na216_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1359_1_i) );
// C_///AND/D      x156y68     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1360_4 ( .OUT(na1360_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1360_5 ( .OUT(na1360_2), .CLK(na2414_1), .EN(na216_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1360_2_i) );
// C_AND/D///      x145y78     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1361_1 ( .OUT(na1361_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1361_2 ( .OUT(na1361_1), .CLK(na2414_1), .EN(na216_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1361_1_i) );
// C_///AND/D      x142y41     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1362_4 ( .OUT(na1362_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1362_5 ( .OUT(na1362_2), .CLK(na2414_1), .EN(na217_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1362_2_i) );
// C_AND/D///      x132y36     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1363_1 ( .OUT(na1363_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1363_2 ( .OUT(na1363_1), .CLK(na2414_1), .EN(na217_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1363_1_i) );
// C_AND/D///      x150y45     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1364_1 ( .OUT(na1364_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2403_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1364_2 ( .OUT(na1364_1), .CLK(na2414_1), .EN(na217_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1364_1_i) );
// C_AND/D///      x139y52     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1365_1 ( .OUT(na1365_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1365_2 ( .OUT(na1365_1), .CLK(na2414_1), .EN(na217_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1365_1_i) );
// C_///AND/D      x149y57     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1366_4 ( .OUT(na1366_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1366_5 ( .OUT(na1366_2), .CLK(na2414_1), .EN(na217_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1366_2_i) );
// C_AND/D///      x155y53     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1367_1 ( .OUT(na1367_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1367_2 ( .OUT(na1367_1), .CLK(na2414_1), .EN(na217_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1367_1_i) );
// C_///AND/D      x144y75     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1368_4 ( .OUT(na1368_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1368_5 ( .OUT(na1368_2), .CLK(na2414_1), .EN(na217_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1368_2_i) );
// C_AND/D///      x149y72     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1369_1 ( .OUT(na1369_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1369_2 ( .OUT(na1369_1), .CLK(na2414_1), .EN(na217_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1369_1_i) );
// C_///AND/D      x155y78     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1370_4 ( .OUT(na1370_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1370_5 ( .OUT(na1370_2), .CLK(na2414_1), .EN(na217_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1370_2_i) );
// C_///AND/D      x138y80     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1371_4 ( .OUT(na1371_2_i), .IN1(1'b1), .IN2(na2410_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1371_5 ( .OUT(na1371_2), .CLK(na2414_1), .EN(na217_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1371_2_i) );
// C_///AND/D      x146y42     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1372_4 ( .OUT(na1372_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1372_5 ( .OUT(na1372_2), .CLK(na2414_1), .EN(na218_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1372_2_i) );
// C_AND/D///      x132y37     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1373_1 ( .OUT(na1373_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1373_2 ( .OUT(na1373_1), .CLK(na2414_1), .EN(na218_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1373_1_i) );
// C_///AND/D      x150y56     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1374_4 ( .OUT(na1374_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1374_5 ( .OUT(na1374_2), .CLK(na2414_1), .EN(na218_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1374_2_i) );
// C_AND/D///      x139y51     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1375_1 ( .OUT(na1375_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1375_2 ( .OUT(na1375_1), .CLK(na2414_1), .EN(na218_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1375_1_i) );
// C_///AND/D      x149y56     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1376_4 ( .OUT(na1376_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1376_5 ( .OUT(na1376_2), .CLK(na2414_1), .EN(na218_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1376_2_i) );
// C_AND/D///      x153y56     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1377_1 ( .OUT(na1377_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1377_2 ( .OUT(na1377_1), .CLK(na2414_1), .EN(na218_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1377_1_i) );
// C_AND/D///      x146y68     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1378_1 ( .OUT(na1378_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2407_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1378_2 ( .OUT(na1378_1), .CLK(na2414_1), .EN(na218_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1378_1_i) );
// C_AND/D///      x151y71     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1379_1 ( .OUT(na1379_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1379_2 ( .OUT(na1379_1), .CLK(na2414_1), .EN(na218_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1379_1_i) );
// C_///AND/D      x151y79     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1380_4 ( .OUT(na1380_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1380_5 ( .OUT(na1380_2), .CLK(na2414_1), .EN(na218_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1380_2_i) );
// C_AND/D///      x144y81     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1381_1 ( .OUT(na1381_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1381_2 ( .OUT(na1381_1), .CLK(na2414_1), .EN(na218_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1381_1_i) );
// C_///AND/D      x149y41     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1382_4 ( .OUT(na1382_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1382_5 ( .OUT(na1382_2), .CLK(na2414_1), .EN(na219_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1382_2_i) );
// C_AND/D///      x135y38     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1383_1 ( .OUT(na1383_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1383_2 ( .OUT(na1383_1), .CLK(na2414_1), .EN(na219_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1383_1_i) );
// C_///AND/D      x149y55     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1384_4 ( .OUT(na1384_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1384_5 ( .OUT(na1384_2), .CLK(na2414_1), .EN(na219_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1384_2_i) );
// C_///AND/D      x136y48     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1385_4 ( .OUT(na1385_2_i), .IN1(1'b1), .IN2(na2404_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1385_5 ( .OUT(na1385_2), .CLK(na2414_1), .EN(na219_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1385_2_i) );
// C_///AND/D      x148y51     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1386_4 ( .OUT(na1386_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1386_5 ( .OUT(na1386_2), .CLK(na2414_1), .EN(na219_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1386_2_i) );
// C_AND/D///      x154y55     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1387_1 ( .OUT(na1387_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1387_2 ( .OUT(na1387_1), .CLK(na2414_1), .EN(na219_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1387_1_i) );
// C_///AND/D      x147y77     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1388_4 ( .OUT(na1388_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1388_5 ( .OUT(na1388_2), .CLK(na2414_1), .EN(na219_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1388_2_i) );
// C_AND/D///      x150y72     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1389_1 ( .OUT(na1389_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1389_2 ( .OUT(na1389_1), .CLK(na2414_1), .EN(na219_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1389_1_i) );
// C_///AND/D      x156y80     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1390_4 ( .OUT(na1390_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1390_5 ( .OUT(na1390_2), .CLK(na2414_1), .EN(na219_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1390_2_i) );
// C_AND/D///      x147y84     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1391_1 ( .OUT(na1391_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1391_2 ( .OUT(na1391_1), .CLK(na2414_1), .EN(na219_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1391_1_i) );
// C_AND/D///      x150y40     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1392_1 ( .OUT(na1392_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2401_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1392_2 ( .OUT(na1392_1), .CLK(na2414_1), .EN(na214_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1392_1_i) );
// C_AND/D///      x132y41     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1393_1 ( .OUT(na1393_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1393_2 ( .OUT(na1393_1), .CLK(na2414_1), .EN(na214_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1393_1_i) );
// C_///AND/D      x143y54     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1394_4 ( .OUT(na1394_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1394_5 ( .OUT(na1394_2), .CLK(na2414_1), .EN(na214_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1394_2_i) );
// C_AND/D///      x137y56     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1395_1 ( .OUT(na1395_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1395_2 ( .OUT(na1395_1), .CLK(na2414_1), .EN(na214_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1395_1_i) );
// C_///AND/D      x148y62     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1396_4 ( .OUT(na1396_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1396_5 ( .OUT(na1396_2), .CLK(na2414_1), .EN(na214_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1396_2_i) );
// C_AND/D///      x154y62     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1397_1 ( .OUT(na1397_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1397_2 ( .OUT(na1397_1), .CLK(na2414_1), .EN(na214_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1397_1_i) );
// C_///AND/D      x149y77     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1398_4 ( .OUT(na1398_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1398_5 ( .OUT(na1398_2), .CLK(na2414_1), .EN(na214_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1398_2_i) );
// C_///AND/D      x149y74     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1399_4 ( .OUT(na1399_2_i), .IN1(na2408_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1399_5 ( .OUT(na1399_2), .CLK(na2414_1), .EN(na214_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1399_2_i) );
// C_///AND/D      x155y70     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1400_4 ( .OUT(na1400_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1400_5 ( .OUT(na1400_2), .CLK(na2414_1), .EN(na214_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1400_2_i) );
// C_AND/D///      x144y78     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1401_1 ( .OUT(na1401_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1401_2 ( .OUT(na1401_1), .CLK(na2414_1), .EN(na214_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1401_1_i) );
// C_///AND/D      x114y38     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1402_4 ( .OUT(na1402_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1402_5 ( .OUT(na1402_2), .CLK(na2414_1), .EN(na237_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1402_2_i) );
// C_AND/D///      x114y38     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1403_1 ( .OUT(na1403_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1403_2 ( .OUT(na1403_1), .CLK(na2414_1), .EN(na237_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1403_1_i) );
// C_///AND/D      x108y43     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1404_4 ( .OUT(na1404_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1404_5 ( .OUT(na1404_2), .CLK(na2414_1), .EN(na237_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1404_2_i) );
// C_AND/D///      x108y46     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1405_1 ( .OUT(na1405_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1405_2 ( .OUT(na1405_1), .CLK(na2414_1), .EN(na237_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1405_1_i) );
// C_AND/D///      x105y59     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1406_1 ( .OUT(na1406_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2405_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1406_2 ( .OUT(na1406_1), .CLK(na2414_1), .EN(na237_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1406_1_i) );
// C_AND/D///      x117y58     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1407_1 ( .OUT(na1407_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1407_2 ( .OUT(na1407_1), .CLK(na2414_1), .EN(na237_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1407_1_i) );
// C_///AND/D      x108y71     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1408_4 ( .OUT(na1408_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1408_5 ( .OUT(na1408_2), .CLK(na2414_1), .EN(na237_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1408_2_i) );
// C_AND/D///      x106y74     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1409_1 ( .OUT(na1409_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1409_2 ( .OUT(na1409_1), .CLK(na2414_1), .EN(na237_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1409_1_i) );
// C_///AND/D      x116y82     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1410_4 ( .OUT(na1410_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1410_5 ( .OUT(na1410_2), .CLK(na2414_1), .EN(na237_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1410_2_i) );
// C_AND/D///      x123y79     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1411_1 ( .OUT(na1411_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1411_2 ( .OUT(na1411_1), .CLK(na2414_1), .EN(na237_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1411_1_i) );
// C_///AND/D      x111y38     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1412_4 ( .OUT(na1412_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1412_5 ( .OUT(na1412_2), .CLK(na2414_1), .EN(na223_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1412_2_i) );
// C_///AND/D      x109y35     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1413_4 ( .OUT(na1413_2_i), .IN1(na2402_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1413_5 ( .OUT(na1413_2), .CLK(na2414_1), .EN(na223_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1413_2_i) );
// C_///AND/D      x106y38     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1414_4 ( .OUT(na1414_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1414_5 ( .OUT(na1414_2), .CLK(na2414_1), .EN(na223_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1414_2_i) );
// C_AND/D///      x110y42     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1415_1 ( .OUT(na1415_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1415_2 ( .OUT(na1415_1), .CLK(na2414_1), .EN(na223_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1415_1_i) );
// C_///AND/D      x107y59     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1416_4 ( .OUT(na1416_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1416_5 ( .OUT(na1416_2), .CLK(na2414_1), .EN(na223_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1416_2_i) );
// C_AND/D///      x114y61     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1417_1 ( .OUT(na1417_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1417_2 ( .OUT(na1417_1), .CLK(na2414_1), .EN(na223_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1417_1_i) );
// C_///AND/D      x107y66     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1418_4 ( .OUT(na1418_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1418_5 ( .OUT(na1418_2), .CLK(na2414_1), .EN(na223_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1418_2_i) );
// C_AND/D///      x106y72     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1419_1 ( .OUT(na1419_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1419_2 ( .OUT(na1419_1), .CLK(na2414_1), .EN(na223_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1419_1_i) );
// C_AND/D///      x109y84     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1420_1 ( .OUT(na1420_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2409_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1420_2 ( .OUT(na1420_1), .CLK(na2414_1), .EN(na223_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1420_1_i) );
// C_AND/D///      x120y83     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1421_1 ( .OUT(na1421_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1421_2 ( .OUT(na1421_1), .CLK(na2414_1), .EN(na223_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1421_1_i) );
// C_///AND/D      x112y35     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1422_4 ( .OUT(na1422_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1422_5 ( .OUT(na1422_2), .CLK(na2414_1), .EN(na224_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1422_2_i) );
// C_AND/D///      x108y34     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1423_1 ( .OUT(na1423_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1423_2 ( .OUT(na1423_1), .CLK(na2414_1), .EN(na224_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1423_1_i) );
// C_///AND/D      x107y37     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1424_4 ( .OUT(na1424_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1424_5 ( .OUT(na1424_2), .CLK(na2414_1), .EN(na224_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1424_2_i) );
// C_AND/D///      x111y43     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1425_1 ( .OUT(na1425_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1425_2 ( .OUT(na1425_1), .CLK(na2414_1), .EN(na224_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1425_1_i) );
// C_///AND/D      x110y58     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1426_4 ( .OUT(na1426_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1426_5 ( .OUT(na1426_2), .CLK(na2414_1), .EN(na224_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1426_2_i) );
// C_///AND/D      x121y62     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1427_4 ( .OUT(na1427_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2406_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1427_5 ( .OUT(na1427_2), .CLK(na2414_1), .EN(na224_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1427_2_i) );
// C_///AND/D      x112y65     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1428_4 ( .OUT(na1428_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1428_5 ( .OUT(na1428_2), .CLK(na2414_1), .EN(na224_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1428_2_i) );
// C_AND/D///      x107y71     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1429_1 ( .OUT(na1429_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1429_2 ( .OUT(na1429_1), .CLK(na2414_1), .EN(na224_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1429_1_i) );
// C_///AND/D      x108y83     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1430_4 ( .OUT(na1430_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1430_5 ( .OUT(na1430_2), .CLK(na2414_1), .EN(na224_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1430_2_i) );
// C_AND/D///      x119y82     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1431_1 ( .OUT(na1431_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1431_2 ( .OUT(na1431_1), .CLK(na2414_1), .EN(na224_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1431_1_i) );
// C_///AND/D      x116y40     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1432_4 ( .OUT(na1432_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1432_5 ( .OUT(na1432_2), .CLK(na2414_1), .EN(na225_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1432_2_i) );
// C_AND/D///      x110y33     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1433_1 ( .OUT(na1433_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1433_2 ( .OUT(na1433_1), .CLK(na2414_1), .EN(na225_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1433_1_i) );
// C_AND/D///      x105y40     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1434_1 ( .OUT(na1434_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2403_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1434_2 ( .OUT(na1434_1), .CLK(na2414_1), .EN(na225_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1434_1_i) );
// C_AND/D///      x109y44     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1435_1 ( .OUT(na1435_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1435_2 ( .OUT(na1435_1), .CLK(na2414_1), .EN(na225_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1435_1_i) );
// C_///AND/D      x110y57     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1436_4 ( .OUT(na1436_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1436_5 ( .OUT(na1436_2), .CLK(na2414_1), .EN(na225_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1436_2_i) );
// C_AND/D///      x113y63     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1437_1 ( .OUT(na1437_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1437_2 ( .OUT(na1437_1), .CLK(na2414_1), .EN(na225_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1437_1_i) );
// C_///AND/D      x108y68     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1438_4 ( .OUT(na1438_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1438_5 ( .OUT(na1438_2), .CLK(na2414_1), .EN(na225_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1438_2_i) );
// C_AND/D///      x107y70     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1439_1 ( .OUT(na1439_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1439_2 ( .OUT(na1439_1), .CLK(na2414_1), .EN(na225_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1439_1_i) );
// C_///AND/D      x108y82     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1440_4 ( .OUT(na1440_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1440_5 ( .OUT(na1440_2), .CLK(na2414_1), .EN(na225_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1440_2_i) );
// C_///AND/D      x129y81     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1441_4 ( .OUT(na1441_2_i), .IN1(1'b1), .IN2(na2410_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1441_5 ( .OUT(na1441_2), .CLK(na2414_1), .EN(na225_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1441_2_i) );
// C_///AND/D      x111y36     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1442_4 ( .OUT(na1442_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1442_5 ( .OUT(na1442_2), .CLK(na2414_1), .EN(na226_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1442_2_i) );
// C_AND/D///      x111y36     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1443_1 ( .OUT(na1443_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1443_2 ( .OUT(na1443_1), .CLK(na2414_1), .EN(na226_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1443_1_i) );
// C_///AND/D      x113y38     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1444_4 ( .OUT(na1444_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1444_5 ( .OUT(na1444_2), .CLK(na2414_1), .EN(na226_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1444_2_i) );
// C_AND/D///      x110y48     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1445_1 ( .OUT(na1445_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1445_2 ( .OUT(na1445_1), .CLK(na2414_1), .EN(na226_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1445_1_i) );
// C_///AND/D      x106y59     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1446_4 ( .OUT(na1446_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1446_5 ( .OUT(na1446_2), .CLK(na2414_1), .EN(na226_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1446_2_i) );
// C_AND/D///      x119y61     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1447_1 ( .OUT(na1447_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1447_2 ( .OUT(na1447_1), .CLK(na2414_1), .EN(na226_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1447_1_i) );
// C_AND/D///      x106y65     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1448_1 ( .OUT(na1448_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2407_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1448_2 ( .OUT(na1448_1), .CLK(na2414_1), .EN(na226_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1448_1_i) );
// C_AND/D///      x105y71     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1449_1 ( .OUT(na1449_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1449_2 ( .OUT(na1449_1), .CLK(na2414_1), .EN(na226_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1449_1_i) );
// C_///AND/D      x116y81     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1450_4 ( .OUT(na1450_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1450_5 ( .OUT(na1450_2), .CLK(na2414_1), .EN(na226_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1450_2_i) );
// C_AND/D///      x121y74     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1451_1 ( .OUT(na1451_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1451_2 ( .OUT(na1451_1), .CLK(na2414_1), .EN(na226_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1451_1_i) );
// C_///AND/D      x111y39     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1452_4 ( .OUT(na1452_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1452_5 ( .OUT(na1452_2), .CLK(na2414_1), .EN(na227_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1452_2_i) );
// C_AND/D///      x111y37     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1453_1 ( .OUT(na1453_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1453_2 ( .OUT(na1453_1), .CLK(na2414_1), .EN(na227_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1453_1_i) );
// C_///AND/D      x107y39     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1454_4 ( .OUT(na1454_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1454_5 ( .OUT(na1454_2), .CLK(na2414_1), .EN(na227_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1454_2_i) );
// C_///AND/D      x114y49     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1455_4 ( .OUT(na1455_2_i), .IN1(1'b1), .IN2(na2404_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1455_5 ( .OUT(na1455_2), .CLK(na2414_1), .EN(na227_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1455_2_i) );
// C_///AND/D      x112y60     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1456_4 ( .OUT(na1456_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1456_5 ( .OUT(na1456_2), .CLK(na2414_1), .EN(na227_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1456_2_i) );
// C_AND/D///      x117y64     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1457_1 ( .OUT(na1457_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1457_2 ( .OUT(na1457_1), .CLK(na2414_1), .EN(na227_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1457_1_i) );
// C_///AND/D      x106y70     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1458_4 ( .OUT(na1458_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1458_5 ( .OUT(na1458_2), .CLK(na2414_1), .EN(na227_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1458_2_i) );
// C_AND/D///      x109y72     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1459_1 ( .OUT(na1459_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1459_2 ( .OUT(na1459_1), .CLK(na2414_1), .EN(na227_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1459_1_i) );
// C_///AND/D      x112y82     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1460_4 ( .OUT(na1460_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1460_5 ( .OUT(na1460_2), .CLK(na2414_1), .EN(na227_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1460_2_i) );
// C_AND/D///      x121y75     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1461_1 ( .OUT(na1461_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1461_2 ( .OUT(na1461_1), .CLK(na2414_1), .EN(na227_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1461_1_i) );
// C_AND/D///      x112y32     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1462_1 ( .OUT(na1462_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2401_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1462_2 ( .OUT(na1462_1), .CLK(na2414_1), .EN(na228_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1462_1_i) );
// C_AND/D///      x112y38     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1463_1 ( .OUT(na1463_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1463_2 ( .OUT(na1463_1), .CLK(na2414_1), .EN(na228_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1463_1_i) );
// C_///AND/D      x108y42     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1464_4 ( .OUT(na1464_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1464_5 ( .OUT(na1464_2), .CLK(na2414_1), .EN(na228_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1464_2_i) );
// C_AND/D///      x111y48     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1465_1 ( .OUT(na1465_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1465_2 ( .OUT(na1465_1), .CLK(na2414_1), .EN(na228_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1465_1_i) );
// C_///AND/D      x107y63     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1466_4 ( .OUT(na1466_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1466_5 ( .OUT(na1466_2), .CLK(na2414_1), .EN(na228_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1466_2_i) );
// C_AND/D///      x120y63     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1467_1 ( .OUT(na1467_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1467_2 ( .OUT(na1467_1), .CLK(na2414_1), .EN(na228_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1467_1_i) );
// C_///AND/D      x107y69     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1468_4 ( .OUT(na1468_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1468_5 ( .OUT(na1468_2), .CLK(na2414_1), .EN(na228_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1468_2_i) );
// C_///AND/D      x112y79     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1469_4 ( .OUT(na1469_2_i), .IN1(na2408_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1469_5 ( .OUT(na1469_2), .CLK(na2414_1), .EN(na228_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1469_2_i) );
// C_///AND/D      x113y81     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1470_4 ( .OUT(na1470_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1470_5 ( .OUT(na1470_2), .CLK(na2414_1), .EN(na228_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1470_2_i) );
// C_AND/D///      x122y76     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1471_1 ( .OUT(na1471_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1471_2 ( .OUT(na1471_1), .CLK(na2414_1), .EN(na228_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1471_1_i) );
// C_///AND/D      x114y39     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1472_4 ( .OUT(na1472_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1472_5 ( .OUT(na1472_2), .CLK(na2414_1), .EN(na229_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1472_2_i) );
// C_AND/D///      x116y37     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1473_1 ( .OUT(na1473_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1473_2 ( .OUT(na1473_1), .CLK(na2414_1), .EN(na229_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1473_1_i) );
// C_///AND/D      x108y39     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1474_4 ( .OUT(na1474_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1474_5 ( .OUT(na1474_2), .CLK(na2414_1), .EN(na229_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1474_2_i) );
// C_AND/D///      x111y47     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1475_1 ( .OUT(na1475_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1475_2 ( .OUT(na1475_1), .CLK(na2414_1), .EN(na229_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1475_1_i) );
// C_AND/D///      x105y60     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1476_1 ( .OUT(na1476_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2405_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1476_2 ( .OUT(na1476_1), .CLK(na2414_1), .EN(na229_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1476_1_i) );
// C_AND/D///      x120y64     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1477_1 ( .OUT(na1477_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1477_2 ( .OUT(na1477_1), .CLK(na2414_1), .EN(na229_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1477_1_i) );
// C_///AND/D      x107y72     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1478_4 ( .OUT(na1478_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1478_5 ( .OUT(na1478_2), .CLK(na2414_1), .EN(na229_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1478_2_i) );
// C_AND/D///      x108y72     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1479_1 ( .OUT(na1479_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1479_2 ( .OUT(na1479_1), .CLK(na2414_1), .EN(na229_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1479_1_i) );
// C_///AND/D      x113y84     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1480_4 ( .OUT(na1480_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1480_5 ( .OUT(na1480_2), .CLK(na2414_1), .EN(na229_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1480_2_i) );
// C_AND/D///      x124y75     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1481_1 ( .OUT(na1481_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1481_2 ( .OUT(na1481_1), .CLK(na2414_1), .EN(na229_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1481_1_i) );
// C_///AND/D      x116y36     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1482_4 ( .OUT(na1482_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1482_5 ( .OUT(na1482_2), .CLK(na2414_1), .EN(na230_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1482_2_i) );
// C_///AND/D      x118y40     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1483_4 ( .OUT(na1483_2_i), .IN1(na2402_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1483_5 ( .OUT(na1483_2), .CLK(na2414_1), .EN(na230_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1483_2_i) );
// C_///AND/D      x111y41     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1484_4 ( .OUT(na1484_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1484_5 ( .OUT(na1484_2), .CLK(na2414_1), .EN(na230_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1484_2_i) );
// C_AND/D///      x111y41     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1485_1 ( .OUT(na1485_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1485_2 ( .OUT(na1485_1), .CLK(na2414_1), .EN(na230_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1485_1_i) );
// C_///AND/D      x110y62     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1486_4 ( .OUT(na1486_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1486_5 ( .OUT(na1486_2), .CLK(na2414_1), .EN(na230_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1486_2_i) );
// C_AND/D///      x114y58     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1487_1 ( .OUT(na1487_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1487_2 ( .OUT(na1487_1), .CLK(na2414_1), .EN(na230_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1487_1_i) );
// C_///AND/D      x112y71     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1488_4 ( .OUT(na1488_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1488_5 ( .OUT(na1488_2), .CLK(na2414_1), .EN(na230_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1488_2_i) );
// C_AND/D///      x107y74     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1489_1 ( .OUT(na1489_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1489_2 ( .OUT(na1489_1), .CLK(na2414_1), .EN(na230_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1489_1_i) );
// C_AND/D///      x114y81     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1490_1 ( .OUT(na1490_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2409_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1490_2 ( .OUT(na1490_1), .CLK(na2414_1), .EN(na230_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1490_1_i) );
// C_AND/D///      x122y80     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1491_1 ( .OUT(na1491_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1491_2 ( .OUT(na1491_1), .CLK(na2414_1), .EN(na230_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1491_1_i) );
// C_///AND/D      x109y39     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1492_4 ( .OUT(na1492_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1492_5 ( .OUT(na1492_2), .CLK(na2414_1), .EN(na221_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1492_2_i) );
// C_AND/D///      x107y34     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1493_1 ( .OUT(na1493_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1493_2 ( .OUT(na1493_1), .CLK(na2414_1), .EN(na221_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1493_1_i) );
// C_///AND/D      x106y39     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1494_4 ( .OUT(na1494_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1494_5 ( .OUT(na1494_2), .CLK(na2414_1), .EN(na221_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1494_2_i) );
// C_AND/D///      x110y43     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1495_1 ( .OUT(na1495_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1495_2 ( .OUT(na1495_1), .CLK(na2414_1), .EN(na221_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1495_1_i) );
// C_///AND/D      x107y62     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1496_4 ( .OUT(na1496_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1496_5 ( .OUT(na1496_2), .CLK(na2414_1), .EN(na221_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1496_2_i) );
// C_///AND/D      x118y64     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1497_4 ( .OUT(na1497_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2406_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1497_5 ( .OUT(na1497_2), .CLK(na2414_1), .EN(na221_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1497_2_i) );
// C_///AND/D      x109y67     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1498_4 ( .OUT(na1498_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1498_5 ( .OUT(na1498_2), .CLK(na2414_1), .EN(na221_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1498_2_i) );
// C_AND/D///      x110y69     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1499_1 ( .OUT(na1499_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1499_2 ( .OUT(na1499_1), .CLK(na2414_1), .EN(na221_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1499_1_i) );
// C_///AND/D      x109y81     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1500_4 ( .OUT(na1500_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1500_5 ( .OUT(na1500_2), .CLK(na2414_1), .EN(na221_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1500_2_i) );
// C_AND/D///      x120y82     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1501_1 ( .OUT(na1501_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1501_2 ( .OUT(na1501_1), .CLK(na2414_1), .EN(na221_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1501_1_i) );
// C_///AND/D      x117y38     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1502_4 ( .OUT(na1502_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1502_5 ( .OUT(na1502_2), .CLK(na2414_1), .EN(na232_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1502_2_i) );
// C_AND/D///      x113y36     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1503_1 ( .OUT(na1503_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1503_2 ( .OUT(na1503_1), .CLK(na2414_1), .EN(na232_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1503_1_i) );
// C_AND/D///      x108y41     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1504_1 ( .OUT(na1504_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2403_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1504_2 ( .OUT(na1504_1), .CLK(na2414_1), .EN(na232_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1504_1_i) );
// C_AND/D///      x112y41     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1505_1 ( .OUT(na1505_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1505_2 ( .OUT(na1505_1), .CLK(na2414_1), .EN(na232_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1505_1_i) );
// C_///AND/D      x113y60     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1506_4 ( .OUT(na1506_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1506_5 ( .OUT(na1506_2), .CLK(na2414_1), .EN(na232_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1506_2_i) );
// C_AND/D///      x115y60     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1507_1 ( .OUT(na1507_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1507_2 ( .OUT(na1507_1), .CLK(na2414_1), .EN(na232_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1507_1_i) );
// C_///AND/D      x109y69     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1508_4 ( .OUT(na1508_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1508_5 ( .OUT(na1508_2), .CLK(na2414_1), .EN(na232_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1508_2_i) );
// C_AND/D///      x108y74     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1509_1 ( .OUT(na1509_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1509_2 ( .OUT(na1509_1), .CLK(na2414_1), .EN(na232_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1509_1_i) );
// C_///AND/D      x119y81     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1510_4 ( .OUT(na1510_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1510_5 ( .OUT(na1510_2), .CLK(na2414_1), .EN(na232_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1510_2_i) );
// C_///AND/D      x123y80     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1511_4 ( .OUT(na1511_2_i), .IN1(1'b1), .IN2(na2410_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1511_5 ( .OUT(na1511_2), .CLK(na2414_1), .EN(na232_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1511_2_i) );
// C_///AND/D      x119y37     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1512_4 ( .OUT(na1512_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1512_5 ( .OUT(na1512_2), .CLK(na2414_1), .EN(na233_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1512_2_i) );
// C_AND/D///      x115y35     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1513_1 ( .OUT(na1513_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1513_2 ( .OUT(na1513_1), .CLK(na2414_1), .EN(na233_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1513_1_i) );
// C_///AND/D      x110y44     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1514_4 ( .OUT(na1514_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1514_5 ( .OUT(na1514_2), .CLK(na2414_1), .EN(na233_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1514_2_i) );
// C_AND/D///      x112y44     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1515_1 ( .OUT(na1515_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1515_2 ( .OUT(na1515_1), .CLK(na2414_1), .EN(na233_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1515_1_i) );
// C_///AND/D      x113y61     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1516_4 ( .OUT(na1516_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1516_5 ( .OUT(na1516_2), .CLK(na2414_1), .EN(na233_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1516_2_i) );
// C_AND/D///      x119y59     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1517_1 ( .OUT(na1517_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1517_2 ( .OUT(na1517_1), .CLK(na2414_1), .EN(na233_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1517_1_i) );
// C_AND/D///      x109y66     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1518_1 ( .OUT(na1518_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2407_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1518_2 ( .OUT(na1518_1), .CLK(na2414_1), .EN(na233_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1518_1_i) );
// C_AND/D///      x110y73     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1519_1 ( .OUT(na1519_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1519_2 ( .OUT(na1519_1), .CLK(na2414_1), .EN(na233_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1519_1_i) );
// C_///AND/D      x119y84     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1520_4 ( .OUT(na1520_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1520_5 ( .OUT(na1520_2), .CLK(na2414_1), .EN(na233_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1520_2_i) );
// C_AND/D///      x121y79     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1521_1 ( .OUT(na1521_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1521_2 ( .OUT(na1521_1), .CLK(na2414_1), .EN(na233_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1521_1_i) );
// C_///AND/D      x121y39     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1522_4 ( .OUT(na1522_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1522_5 ( .OUT(na1522_2), .CLK(na2414_1), .EN(na234_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1522_2_i) );
// C_AND/D///      x115y39     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1523_1 ( .OUT(na1523_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1523_2 ( .OUT(na1523_1), .CLK(na2414_1), .EN(na234_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1523_1_i) );
// C_///AND/D      x105y42     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1524_4 ( .OUT(na1524_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1524_5 ( .OUT(na1524_2), .CLK(na2414_1), .EN(na234_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1524_2_i) );
// C_///AND/D      x109y49     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1525_4 ( .OUT(na1525_2_i), .IN1(1'b1), .IN2(na2404_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1525_5 ( .OUT(na1525_2), .CLK(na2414_1), .EN(na234_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1525_2_i) );
// C_///AND/D      x108y64     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1526_4 ( .OUT(na1526_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1526_5 ( .OUT(na1526_2), .CLK(na2414_1), .EN(na234_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1526_2_i) );
// C_AND/D///      x118y59     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1527_1 ( .OUT(na1527_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1527_2 ( .OUT(na1527_1), .CLK(na2414_1), .EN(na234_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1527_1_i) );
// C_///AND/D      x109y70     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1528_4 ( .OUT(na1528_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1528_5 ( .OUT(na1528_2), .CLK(na2414_1), .EN(na234_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1528_2_i) );
// C_AND/D///      x105y75     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1529_1 ( .OUT(na1529_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1529_2 ( .OUT(na1529_1), .CLK(na2414_1), .EN(na234_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1529_1_i) );
// C_///AND/D      x117y81     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1530_4 ( .OUT(na1530_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1530_5 ( .OUT(na1530_2), .CLK(na2414_1), .EN(na234_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1530_2_i) );
// C_AND/D///      x126y80     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1531_1 ( .OUT(na1531_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1531_2 ( .OUT(na1531_1), .CLK(na2414_1), .EN(na234_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1531_1_i) );
// C_AND/D///      x117y32     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1532_1 ( .OUT(na1532_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2401_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1532_2 ( .OUT(na1532_1), .CLK(na2414_1), .EN(na235_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1532_1_i) );
// C_AND/D///      x115y40     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1533_1 ( .OUT(na1533_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1533_2 ( .OUT(na1533_1), .CLK(na2414_1), .EN(na235_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1533_1_i) );
// C_///AND/D      x107y43     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1534_4 ( .OUT(na1534_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1534_5 ( .OUT(na1534_2), .CLK(na2414_1), .EN(na235_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1534_2_i) );
// C_AND/D///      x109y46     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1535_1 ( .OUT(na1535_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1535_2 ( .OUT(na1535_1), .CLK(na2414_1), .EN(na235_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1535_1_i) );
// C_///AND/D      x112y61     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1536_4 ( .OUT(na1536_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1536_5 ( .OUT(na1536_2), .CLK(na2414_1), .EN(na235_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1536_2_i) );
// C_AND/D///      x118y58     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1537_1 ( .OUT(na1537_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1537_2 ( .OUT(na1537_1), .CLK(na2414_1), .EN(na235_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1537_1_i) );
// C_///AND/D      x107y73     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1538_4 ( .OUT(na1538_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1538_5 ( .OUT(na1538_2), .CLK(na2414_1), .EN(na235_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1538_2_i) );
// C_///AND/D      x109y80     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1539_4 ( .OUT(na1539_2_i), .IN1(na2408_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1539_5 ( .OUT(na1539_2), .CLK(na2414_1), .EN(na235_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1539_2_i) );
// C_///AND/D      x117y82     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1540_4 ( .OUT(na1540_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1540_5 ( .OUT(na1540_2), .CLK(na2414_1), .EN(na235_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1540_2_i) );
// C_AND/D///      x124y79     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1541_1 ( .OUT(na1541_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1541_2 ( .OUT(na1541_1), .CLK(na2414_1), .EN(na235_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1541_1_i) );
// C_///AND/D      x118y41     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1542_4 ( .OUT(na1542_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1542_5 ( .OUT(na1542_2), .CLK(na2414_1), .EN(na236_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1542_2_i) );
// C_AND/D///      x116y39     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1543_1 ( .OUT(na1543_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1543_2 ( .OUT(na1543_1), .CLK(na2414_1), .EN(na236_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1543_1_i) );
// C_///AND/D      x106y44     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1544_4 ( .OUT(na1544_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1544_5 ( .OUT(na1544_2), .CLK(na2414_1), .EN(na236_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1544_2_i) );
// C_AND/D///      x108y47     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1545_1 ( .OUT(na1545_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1545_2 ( .OUT(na1545_1), .CLK(na2414_1), .EN(na236_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1545_1_i) );
// C_AND/D///      x109y60     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1546_1 ( .OUT(na1546_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2405_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1546_2 ( .OUT(na1546_1), .CLK(na2414_1), .EN(na236_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1546_1_i) );
// C_AND/D///      x119y63     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1547_1 ( .OUT(na1547_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1547_2 ( .OUT(na1547_1), .CLK(na2414_1), .EN(na236_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1547_1_i) );
// C_///AND/D      x104y74     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1548_4 ( .OUT(na1548_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1548_5 ( .OUT(na1548_2), .CLK(na2414_1), .EN(na236_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1548_2_i) );
// C_AND/D///      x110y75     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1549_1 ( .OUT(na1549_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1549_2 ( .OUT(na1549_1), .CLK(na2414_1), .EN(na236_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1549_1_i) );
// C_///AND/D      x122y83     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1550_4 ( .OUT(na1550_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1550_5 ( .OUT(na1550_2), .CLK(na2414_1), .EN(na236_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1550_2_i) );
// C_AND/D///      x125y80     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1551_1 ( .OUT(na1551_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1551_2 ( .OUT(na1551_1), .CLK(na2414_1), .EN(na236_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1551_1_i) );
// C_///AND/D      x124y39     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1552_4 ( .OUT(na1552_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1552_5 ( .OUT(na1552_2), .CLK(na2414_1), .EN(na231_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1552_2_i) );
// C_///AND/D      x114y41     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1553_4 ( .OUT(na1553_2_i), .IN1(na2402_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1553_5 ( .OUT(na1553_2), .CLK(na2414_1), .EN(na231_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1553_2_i) );
// C_///AND/D      x107y46     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1554_4 ( .OUT(na1554_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1554_5 ( .OUT(na1554_2), .CLK(na2414_1), .EN(na231_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1554_2_i) );
// C_AND/D///      x111y46     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1555_1 ( .OUT(na1555_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1555_2 ( .OUT(na1555_1), .CLK(na2414_1), .EN(na231_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1555_1_i) );
// C_///AND/D      x108y59     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1556_4 ( .OUT(na1556_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1556_5 ( .OUT(na1556_2), .CLK(na2414_1), .EN(na231_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1556_2_i) );
// C_AND/D///      x116y61     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1557_1 ( .OUT(na1557_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1557_2 ( .OUT(na1557_1), .CLK(na2414_1), .EN(na231_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1557_1_i) );
// C_///AND/D      x112y76     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1558_4 ( .OUT(na1558_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1558_5 ( .OUT(na1558_2), .CLK(na2414_1), .EN(na231_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1558_2_i) );
// C_AND/D///      x111y75     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1559_1 ( .OUT(na1559_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1559_2 ( .OUT(na1559_1), .CLK(na2414_1), .EN(na231_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1559_1_i) );
// C_AND/D///      x114y82     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1560_1 ( .OUT(na1560_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2409_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1560_2 ( .OUT(na1560_1), .CLK(na2414_1), .EN(na231_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1560_1_i) );
// C_AND/D///      x122y77     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1561_1 ( .OUT(na1561_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1561_2 ( .OUT(na1561_1), .CLK(na2414_1), .EN(na231_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1561_1_i) );
// C_///AND/D      x151y31     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1562_4 ( .OUT(na1562_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1562_5 ( .OUT(na1562_2), .CLK(na2414_1), .EN(na254_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1562_2_i) );
// C_AND/D///      x132y34     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1563_1 ( .OUT(na1563_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1563_2 ( .OUT(na1563_1), .CLK(na2414_1), .EN(na254_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1563_1_i) );
// C_///AND/D      x130y42     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1564_4 ( .OUT(na1564_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1564_5 ( .OUT(na1564_2), .CLK(na2414_1), .EN(na254_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1564_2_i) );
// C_AND/D///      x137y47     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1565_1 ( .OUT(na1565_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1565_2 ( .OUT(na1565_1), .CLK(na2414_1), .EN(na254_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1565_1_i) );
// C_///AND/D      x139y65     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1566_4 ( .OUT(na1566_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1566_5 ( .OUT(na1566_2), .CLK(na2414_1), .EN(na254_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1566_2_i) );
// C_///AND/D      x133y64     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1567_4 ( .OUT(na1567_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2406_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1567_5 ( .OUT(na1567_2), .CLK(na2414_1), .EN(na254_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1567_2_i) );
// C_///AND/D      x130y65     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1568_4 ( .OUT(na1568_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1568_5 ( .OUT(na1568_2), .CLK(na2414_1), .EN(na254_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1568_2_i) );
// C_AND/D///      x133y69     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1569_1 ( .OUT(na1569_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1569_2 ( .OUT(na1569_1), .CLK(na2414_1), .EN(na254_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1569_1_i) );
// C_///AND/D      x136y81     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1570_4 ( .OUT(na1570_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1570_5 ( .OUT(na1570_2), .CLK(na2414_1), .EN(na254_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1570_2_i) );
// C_AND/D///      x150y82     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1571_1 ( .OUT(na1571_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1571_2 ( .OUT(na1571_1), .CLK(na2414_1), .EN(na254_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1571_1_i) );
// C_///AND/D      x149y31     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1572_4 ( .OUT(na1572_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1572_5 ( .OUT(na1572_2), .CLK(na2414_1), .EN(na240_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1572_2_i) );
// C_AND/D///      x134y33     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1573_1 ( .OUT(na1573_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1573_2 ( .OUT(na1573_1), .CLK(na2414_1), .EN(na240_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1573_1_i) );
// C_AND/D///      x127y43     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1574_1 ( .OUT(na1574_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2403_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1574_2 ( .OUT(na1574_1), .CLK(na2414_1), .EN(na240_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1574_1_i) );
// C_AND/D///      x138y41     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1575_1 ( .OUT(na1575_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1575_2 ( .OUT(na1575_1), .CLK(na2414_1), .EN(na240_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1575_1_i) );
// C_///AND/D      x129y61     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1576_4 ( .OUT(na1576_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1576_5 ( .OUT(na1576_2), .CLK(na2414_1), .EN(na240_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1576_2_i) );
// C_AND/D///      x135y60     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1577_1 ( .OUT(na1577_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1577_2 ( .OUT(na1577_1), .CLK(na2414_1), .EN(na240_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1577_1_i) );
// C_///AND/D      x128y78     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1578_4 ( .OUT(na1578_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1578_5 ( .OUT(na1578_2), .CLK(na2414_1), .EN(na240_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1578_2_i) );
// C_AND/D///      x128y67     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1579_1 ( .OUT(na1579_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1579_2 ( .OUT(na1579_1), .CLK(na2414_1), .EN(na240_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1579_1_i) );
// C_///AND/D      x133y79     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1580_4 ( .OUT(na1580_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1580_5 ( .OUT(na1580_2), .CLK(na2414_1), .EN(na240_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1580_2_i) );
// C_///AND/D      x141y82     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1581_4 ( .OUT(na1581_2_i), .IN1(1'b1), .IN2(na2410_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1581_5 ( .OUT(na1581_2), .CLK(na2414_1), .EN(na240_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1581_2_i) );
// C_///AND/D      x152y30     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1582_4 ( .OUT(na1582_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1582_5 ( .OUT(na1582_2), .CLK(na2414_1), .EN(na241_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1582_2_i) );
// C_AND/D///      x133y36     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1583_1 ( .OUT(na1583_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1583_2 ( .OUT(na1583_1), .CLK(na2414_1), .EN(na241_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1583_1_i) );
// C_///AND/D      x128y46     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1584_4 ( .OUT(na1584_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1584_5 ( .OUT(na1584_2), .CLK(na2414_1), .EN(na241_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1584_2_i) );
// C_AND/D///      x141y42     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1585_1 ( .OUT(na1585_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1585_2 ( .OUT(na1585_1), .CLK(na2414_1), .EN(na241_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1585_1_i) );
// C_///AND/D      x130y62     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1586_4 ( .OUT(na1586_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1586_5 ( .OUT(na1586_2), .CLK(na2414_1), .EN(na241_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1586_2_i) );
// C_AND/D///      x136y59     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1587_1 ( .OUT(na1587_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1587_2 ( .OUT(na1587_1), .CLK(na2414_1), .EN(na241_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1587_1_i) );
// C_AND/D///      x127y69     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1588_1 ( .OUT(na1588_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2407_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1588_2 ( .OUT(na1588_1), .CLK(na2414_1), .EN(na241_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1588_1_i) );
// C_AND/D///      x129y68     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1589_1 ( .OUT(na1589_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1589_2 ( .OUT(na1589_1), .CLK(na2414_1), .EN(na241_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1589_1_i) );
// C_///AND/D      x136y80     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1590_4 ( .OUT(na1590_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1590_5 ( .OUT(na1590_2), .CLK(na2414_1), .EN(na241_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1590_2_i) );
// C_AND/D///      x148y81     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1591_1 ( .OUT(na1591_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1591_2 ( .OUT(na1591_1), .CLK(na2414_1), .EN(na241_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1591_1_i) );
// C_///AND/D      x150y31     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1592_4 ( .OUT(na1592_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1592_5 ( .OUT(na1592_2), .CLK(na2414_1), .EN(na242_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1592_2_i) );
// C_AND/D///      x135y35     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1593_1 ( .OUT(na1593_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1593_2 ( .OUT(na1593_1), .CLK(na2414_1), .EN(na242_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1593_1_i) );
// C_///AND/D      x126y45     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1594_4 ( .OUT(na1594_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1594_5 ( .OUT(na1594_2), .CLK(na2414_1), .EN(na242_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1594_2_i) );
// C_///AND/D      x133y45     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1595_4 ( .OUT(na1595_2_i), .IN1(1'b1), .IN2(na2404_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1595_5 ( .OUT(na1595_2), .CLK(na2414_1), .EN(na242_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1595_2_i) );
// C_///AND/D      x128y63     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1596_4 ( .OUT(na1596_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1596_5 ( .OUT(na1596_2), .CLK(na2414_1), .EN(na242_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1596_2_i) );
// C_AND/D///      x140y56     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1597_1 ( .OUT(na1597_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1597_2 ( .OUT(na1597_1), .CLK(na2414_1), .EN(na242_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1597_1_i) );
// C_///AND/D      x127y76     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1598_4 ( .OUT(na1598_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1598_5 ( .OUT(na1598_2), .CLK(na2414_1), .EN(na242_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1598_2_i) );
// C_AND/D///      x129y67     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1599_1 ( .OUT(na1599_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1599_2 ( .OUT(na1599_1), .CLK(na2414_1), .EN(na242_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1599_1_i) );
// C_///AND/D      x134y79     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1600_4 ( .OUT(na1600_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1600_5 ( .OUT(na1600_2), .CLK(na2414_1), .EN(na242_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1600_2_i) );
// C_AND/D///      x146y82     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1601_1 ( .OUT(na1601_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1601_2 ( .OUT(na1601_1), .CLK(na2414_1), .EN(na242_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1601_1_i) );
// C_AND/D///      x130y31     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1602_1 ( .OUT(na1602_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2401_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1602_2 ( .OUT(na1602_1), .CLK(na2414_1), .EN(na243_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1602_1_i) );
// C_AND/D///      x135y39     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1603_1 ( .OUT(na1603_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1603_2 ( .OUT(na1603_1), .CLK(na2414_1), .EN(na243_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1603_1_i) );
// C_///AND/D      x128y42     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1604_4 ( .OUT(na1604_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1604_5 ( .OUT(na1604_2), .CLK(na2414_1), .EN(na243_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1604_2_i) );
// C_AND/D///      x136y43     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1605_1 ( .OUT(na1605_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1605_2 ( .OUT(na1605_1), .CLK(na2414_1), .EN(na243_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1605_1_i) );
// C_///AND/D      x133y66     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1606_4 ( .OUT(na1606_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1606_5 ( .OUT(na1606_2), .CLK(na2414_1), .EN(na243_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1606_2_i) );
// C_AND/D///      x139y59     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1607_1 ( .OUT(na1607_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1607_2 ( .OUT(na1607_1), .CLK(na2414_1), .EN(na243_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1607_1_i) );
// C_///AND/D      x119y71     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1608_4 ( .OUT(na1608_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1608_5 ( .OUT(na1608_2), .CLK(na2414_1), .EN(na243_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1608_2_i) );
// C_///AND/D      x138y69     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1609_4 ( .OUT(na1609_2_i), .IN1(na2408_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1609_5 ( .OUT(na1609_2), .CLK(na2414_1), .EN(na243_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1609_2_i) );
// C_///AND/D      x139y79     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1610_4 ( .OUT(na1610_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1610_5 ( .OUT(na1610_2), .CLK(na2414_1), .EN(na243_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1610_2_i) );
// C_AND/D///      x141y81     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1611_1 ( .OUT(na1611_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1611_2 ( .OUT(na1611_1), .CLK(na2414_1), .EN(na243_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1611_1_i) );
// C_///AND/D      x144y32     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1612_4 ( .OUT(na1612_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1612_5 ( .OUT(na1612_2), .CLK(na2414_1), .EN(na244_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1612_2_i) );
// C_AND/D///      x135y40     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1613_1 ( .OUT(na1613_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1613_2 ( .OUT(na1613_1), .CLK(na2414_1), .EN(na244_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1613_1_i) );
// C_///AND/D      x124y43     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1614_4 ( .OUT(na1614_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1614_5 ( .OUT(na1614_2), .CLK(na2414_1), .EN(na244_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1614_2_i) );
// C_AND/D///      x138y46     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1615_1 ( .OUT(na1615_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1615_2 ( .OUT(na1615_1), .CLK(na2414_1), .EN(na244_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1615_1_i) );
// C_AND/D///      x127y63     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1616_1 ( .OUT(na1616_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2405_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1616_2 ( .OUT(na1616_1), .CLK(na2414_1), .EN(na244_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1616_1_i) );
// C_AND/D///      x139y60     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1617_1 ( .OUT(na1617_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1617_2 ( .OUT(na1617_1), .CLK(na2414_1), .EN(na244_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1617_1_i) );
// C_///AND/D      x127y70     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1618_4 ( .OUT(na1618_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1618_5 ( .OUT(na1618_2), .CLK(na2414_1), .EN(na244_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1618_2_i) );
// C_AND/D///      x132y68     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1619_1 ( .OUT(na1619_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1619_2 ( .OUT(na1619_1), .CLK(na2414_1), .EN(na244_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1619_1_i) );
// C_///AND/D      x141y78     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1620_4 ( .OUT(na1620_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1620_5 ( .OUT(na1620_2), .CLK(na2414_1), .EN(na244_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1620_2_i) );
// C_AND/D///      x139y82     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1621_1 ( .OUT(na1621_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1621_2 ( .OUT(na1621_1), .CLK(na2414_1), .EN(na244_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1621_1_i) );
// C_///AND/D      x147y31     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1622_4 ( .OUT(na1622_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1622_5 ( .OUT(na1622_2), .CLK(na2414_1), .EN(na245_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1622_2_i) );
// C_///AND/D      x126y37     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1623_4 ( .OUT(na1623_2_i), .IN1(na2402_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1623_5 ( .OUT(na1623_2), .CLK(na2414_1), .EN(na245_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1623_2_i) );
// C_///AND/D      x123y40     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1624_4 ( .OUT(na1624_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1624_5 ( .OUT(na1624_2), .CLK(na2414_1), .EN(na245_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1624_2_i) );
// C_AND/D///      x137y43     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1625_1 ( .OUT(na1625_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1625_2 ( .OUT(na1625_1), .CLK(na2414_1), .EN(na245_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1625_1_i) );
// C_///AND/D      x134y66     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1626_4 ( .OUT(na1626_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1626_5 ( .OUT(na1626_2), .CLK(na2414_1), .EN(na245_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1626_2_i) );
// C_AND/D///      x138y61     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1627_1 ( .OUT(na1627_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1627_2 ( .OUT(na1627_1), .CLK(na2414_1), .EN(na245_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1627_1_i) );
// C_///AND/D      x132y71     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1628_4 ( .OUT(na1628_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1628_5 ( .OUT(na1628_2), .CLK(na2414_1), .EN(na245_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1628_2_i) );
// C_AND/D///      x129y69     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1629_1 ( .OUT(na1629_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1629_2 ( .OUT(na1629_1), .CLK(na2414_1), .EN(na245_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1629_1_i) );
// C_AND/D///      x138y73     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1630_1 ( .OUT(na1630_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2409_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1630_2 ( .OUT(na1630_1), .CLK(na2414_1), .EN(na245_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1630_1_i) );
// C_AND/D///      x144y83     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1631_1 ( .OUT(na1631_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1631_2 ( .OUT(na1631_1), .CLK(na2414_1), .EN(na245_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1631_1_i) );
// C_///AND/D      x133y34     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1632_4 ( .OUT(na1632_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1632_5 ( .OUT(na1632_2), .CLK(na2414_1), .EN(na246_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1632_2_i) );
// C_AND/D///      x138y40     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1633_1 ( .OUT(na1633_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1633_2 ( .OUT(na1633_1), .CLK(na2414_1), .EN(na246_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1633_1_i) );
// C_///AND/D      x125y45     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1634_4 ( .OUT(na1634_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1634_5 ( .OUT(na1634_2), .CLK(na2414_1), .EN(na246_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1634_2_i) );
// C_AND/D///      x139y44     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1635_1 ( .OUT(na1635_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1635_2 ( .OUT(na1635_1), .CLK(na2414_1), .EN(na246_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1635_1_i) );
// C_///AND/D      x132y69     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1636_4 ( .OUT(na1636_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1636_5 ( .OUT(na1636_2), .CLK(na2414_1), .EN(na246_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1636_2_i) );
// C_///AND/D      x132y62     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1637_4 ( .OUT(na1637_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2406_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1637_5 ( .OUT(na1637_2), .CLK(na2414_1), .EN(na246_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1637_2_i) );
// C_///AND/D      x126y74     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1638_4 ( .OUT(na1638_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1638_5 ( .OUT(na1638_2), .CLK(na2414_1), .EN(na246_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1638_2_i) );
// C_AND/D///      x131y70     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1639_1 ( .OUT(na1639_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1639_2 ( .OUT(na1639_1), .CLK(na2414_1), .EN(na246_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1639_1_i) );
// C_///AND/D      x138y78     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1640_4 ( .OUT(na1640_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1640_5 ( .OUT(na1640_2), .CLK(na2414_1), .EN(na246_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1640_2_i) );
// C_AND/D///      x144y82     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1641_1 ( .OUT(na1641_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1641_2 ( .OUT(na1641_1), .CLK(na2414_1), .EN(na246_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1641_1_i) );
// C_///AND/D      x153y31     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1642_4 ( .OUT(na1642_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1642_5 ( .OUT(na1642_2), .CLK(na2414_1), .EN(na247_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1642_2_i) );
// C_AND/D///      x138y34     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1643_1 ( .OUT(na1643_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1643_2 ( .OUT(na1643_1), .CLK(na2414_1), .EN(na247_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1643_1_i) );
// C_AND/D///      x126y40     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1644_1 ( .OUT(na1644_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2403_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1644_2 ( .OUT(na1644_1), .CLK(na2414_1), .EN(na247_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1644_1_i) );
// C_AND/D///      x140y48     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1645_1 ( .OUT(na1645_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1645_2 ( .OUT(na1645_1), .CLK(na2414_1), .EN(na247_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1645_1_i) );
// C_///AND/D      x141y65     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1646_4 ( .OUT(na1646_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1646_5 ( .OUT(na1646_2), .CLK(na2414_1), .EN(na247_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1646_2_i) );
// C_AND/D///      x136y62     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1647_1 ( .OUT(na1647_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1647_2 ( .OUT(na1647_1), .CLK(na2414_1), .EN(na247_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1647_1_i) );
// C_///AND/D      x129y74     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1648_4 ( .OUT(na1648_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1648_5 ( .OUT(na1648_2), .CLK(na2414_1), .EN(na247_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1648_2_i) );
// C_AND/D///      x134y73     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1649_1 ( .OUT(na1649_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1649_2 ( .OUT(na1649_1), .CLK(na2414_1), .EN(na247_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1649_1_i) );
// C_///AND/D      x134y77     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1650_4 ( .OUT(na1650_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1650_5 ( .OUT(na1650_2), .CLK(na2414_1), .EN(na247_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1650_2_i) );
// C_///AND/D      x142y84     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1651_4 ( .OUT(na1651_2_i), .IN1(1'b1), .IN2(na2410_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1651_5 ( .OUT(na1651_2), .CLK(na2414_1), .EN(na247_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1651_2_i) );
// C_///AND/D      x149y34     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1652_4 ( .OUT(na1652_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1652_5 ( .OUT(na1652_2), .CLK(na2414_1), .EN(na238_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1652_2_i) );
// C_AND/D///      x134y36     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1653_1 ( .OUT(na1653_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1653_2 ( .OUT(na1653_1), .CLK(na2414_1), .EN(na238_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1653_1_i) );
// C_///AND/D      x127y48     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1654_4 ( .OUT(na1654_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1654_5 ( .OUT(na1654_2), .CLK(na2414_1), .EN(na238_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1654_2_i) );
// C_AND/D///      x140y42     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1655_1 ( .OUT(na1655_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1655_2 ( .OUT(na1655_1), .CLK(na2414_1), .EN(na238_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1655_1_i) );
// C_///AND/D      x131y64     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1656_4 ( .OUT(na1656_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1656_5 ( .OUT(na1656_2), .CLK(na2414_1), .EN(na238_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1656_2_i) );
// C_AND/D///      x139y57     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1657_1 ( .OUT(na1657_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1657_2 ( .OUT(na1657_1), .CLK(na2414_1), .EN(na238_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1657_1_i) );
// C_AND/D///      x128y71     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1658_1 ( .OUT(na1658_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2407_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1658_2 ( .OUT(na1658_1), .CLK(na2414_1), .EN(na238_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1658_1_i) );
// C_AND/D///      x130y70     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1659_1 ( .OUT(na1659_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1659_2 ( .OUT(na1659_1), .CLK(na2414_1), .EN(na238_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1659_1_i) );
// C_///AND/D      x137y82     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1660_4 ( .OUT(na1660_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1660_5 ( .OUT(na1660_2), .CLK(na2414_1), .EN(na238_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1660_2_i) );
// C_AND/D///      x147y81     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1661_1 ( .OUT(na1661_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1661_2 ( .OUT(na1661_1), .CLK(na2414_1), .EN(na238_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1661_1_i) );
// C_///AND/D      x156y31     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1662_4 ( .OUT(na1662_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1662_5 ( .OUT(na1662_2), .CLK(na2414_1), .EN(na249_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1662_2_i) );
// C_AND/D///      x137y36     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1663_1 ( .OUT(na1663_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1663_2 ( .OUT(na1663_1), .CLK(na2414_1), .EN(na249_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1663_1_i) );
// C_///AND/D      x129y42     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1664_4 ( .OUT(na1664_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1664_5 ( .OUT(na1664_2), .CLK(na2414_1), .EN(na249_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1664_2_i) );
// C_///AND/D      x131y48     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1665_4 ( .OUT(na1665_2_i), .IN1(1'b1), .IN2(na2404_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1665_5 ( .OUT(na1665_2), .CLK(na2414_1), .EN(na249_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1665_2_i) );
// C_///AND/D      x138y65     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1666_4 ( .OUT(na1666_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1666_5 ( .OUT(na1666_2), .CLK(na2414_1), .EN(na249_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1666_2_i) );
// C_AND/D///      x139y62     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1667_1 ( .OUT(na1667_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1667_2 ( .OUT(na1667_1), .CLK(na2414_1), .EN(na249_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1667_1_i) );
// C_///AND/D      x124y80     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1668_4 ( .OUT(na1668_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1668_5 ( .OUT(na1668_2), .CLK(na2414_1), .EN(na249_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1668_2_i) );
// C_AND/D///      x135y71     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1669_1 ( .OUT(na1669_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1669_2 ( .OUT(na1669_1), .CLK(na2414_1), .EN(na249_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1669_1_i) );
// C_///AND/D      x137y79     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1670_4 ( .OUT(na1670_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1670_5 ( .OUT(na1670_2), .CLK(na2414_1), .EN(na249_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1670_2_i) );
// C_AND/D///      x153y82     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1671_1 ( .OUT(na1671_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1671_2 ( .OUT(na1671_1), .CLK(na2414_1), .EN(na249_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1671_1_i) );
// C_AND/D///      x138y32     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1672_1 ( .OUT(na1672_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2401_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1672_2 ( .OUT(na1672_1), .CLK(na2414_1), .EN(na250_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1672_1_i) );
// C_AND/D///      x139y35     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1673_1 ( .OUT(na1673_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1673_2 ( .OUT(na1673_1), .CLK(na2414_1), .EN(na250_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1673_1_i) );
// C_///AND/D      x123y43     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1674_4 ( .OUT(na1674_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1674_5 ( .OUT(na1674_2), .CLK(na2414_1), .EN(na250_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1674_2_i) );
// C_AND/D///      x137y45     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1675_1 ( .OUT(na1675_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1675_2 ( .OUT(na1675_1), .CLK(na2414_1), .EN(na250_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1675_1_i) );
// C_///AND/D      x138y68     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1676_4 ( .OUT(na1676_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1676_5 ( .OUT(na1676_2), .CLK(na2414_1), .EN(na250_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1676_2_i) );
// C_AND/D///      x137y63     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1677_1 ( .OUT(na1677_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1677_2 ( .OUT(na1677_1), .CLK(na2414_1), .EN(na250_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1677_1_i) );
// C_///AND/D      x128y79     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1678_4 ( .OUT(na1678_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1678_5 ( .OUT(na1678_2), .CLK(na2414_1), .EN(na250_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1678_2_i) );
// C_///AND/D      x137y76     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1679_4 ( .OUT(na1679_2_i), .IN1(na2408_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1679_5 ( .OUT(na1679_2), .CLK(na2414_1), .EN(na250_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1679_2_i) );
// C_///AND/D      x137y78     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1680_4 ( .OUT(na1680_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1680_5 ( .OUT(na1680_2), .CLK(na2414_1), .EN(na250_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1680_2_i) );
// C_AND/D///      x155y81     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1681_1 ( .OUT(na1681_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1681_2 ( .OUT(na1681_1), .CLK(na2414_1), .EN(na250_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1681_1_i) );
// C_///AND/D      x138y36     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1682_4 ( .OUT(na1682_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1682_5 ( .OUT(na1682_2), .CLK(na2414_1), .EN(na251_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1682_2_i) );
// C_AND/D///      x135y33     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1683_1 ( .OUT(na1683_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1683_2 ( .OUT(na1683_1), .CLK(na2414_1), .EN(na251_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1683_1_i) );
// C_///AND/D      x129y43     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1684_4 ( .OUT(na1684_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1684_5 ( .OUT(na1684_2), .CLK(na2414_1), .EN(na251_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1684_2_i) );
// C_AND/D///      x140y50     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1685_1 ( .OUT(na1685_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1685_2 ( .OUT(na1685_1), .CLK(na2414_1), .EN(na251_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1685_1_i) );
// C_AND/D///      x132y64     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1686_1 ( .OUT(na1686_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2405_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1686_2 ( .OUT(na1686_1), .CLK(na2414_1), .EN(na251_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1686_1_i) );
// C_AND/D///      x140y63     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1687_1 ( .OUT(na1687_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1687_2 ( .OUT(na1687_1), .CLK(na2414_1), .EN(na251_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1687_1_i) );
// C_///AND/D      x127y68     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1688_4 ( .OUT(na1688_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1688_5 ( .OUT(na1688_2), .CLK(na2414_1), .EN(na251_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1688_2_i) );
// C_AND/D///      x138y70     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1689_1 ( .OUT(na1689_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1689_2 ( .OUT(na1689_1), .CLK(na2414_1), .EN(na251_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1689_1_i) );
// C_///AND/D      x133y84     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1690_4 ( .OUT(na1690_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1690_5 ( .OUT(na1690_2), .CLK(na2414_1), .EN(na251_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1690_2_i) );
// C_AND/D///      x151y81     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1691_1 ( .OUT(na1691_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1691_2 ( .OUT(na1691_1), .CLK(na2414_1), .EN(na251_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1691_1_i) );
// C_///AND/D      x136y33     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1692_4 ( .OUT(na1692_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1692_5 ( .OUT(na1692_2), .CLK(na2414_1), .EN(na252_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1692_2_i) );
// C_///AND/D      x133y40     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1693_4 ( .OUT(na1693_2_i), .IN1(na2402_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1693_5 ( .OUT(na1693_2), .CLK(na2414_1), .EN(na252_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1693_2_i) );
// C_///AND/D      x131y44     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1694_4 ( .OUT(na1694_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1694_5 ( .OUT(na1694_2), .CLK(na2414_1), .EN(na252_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1694_2_i) );
// C_AND/D///      x140y49     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1695_1 ( .OUT(na1695_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1695_2 ( .OUT(na1695_1), .CLK(na2414_1), .EN(na252_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1695_1_i) );
// C_///AND/D      x138y67     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1696_4 ( .OUT(na1696_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1696_5 ( .OUT(na1696_2), .CLK(na2414_1), .EN(na252_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1696_2_i) );
// C_AND/D///      x140y64     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1697_1 ( .OUT(na1697_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1697_2 ( .OUT(na1697_1), .CLK(na2414_1), .EN(na252_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1697_1_i) );
// C_///AND/D      x131y67     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1698_4 ( .OUT(na1698_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1698_5 ( .OUT(na1698_2), .CLK(na2414_1), .EN(na252_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1698_2_i) );
// C_AND/D///      x134y69     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1699_1 ( .OUT(na1699_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1699_2 ( .OUT(na1699_1), .CLK(na2414_1), .EN(na252_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1699_1_i) );
// C_AND/D///      x135y75     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1700_1 ( .OUT(na1700_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2409_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1700_2 ( .OUT(na1700_1), .CLK(na2414_1), .EN(na252_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1700_1_i) );
// C_AND/D///      x149y82     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1701_1 ( .OUT(na1701_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1701_2 ( .OUT(na1701_1), .CLK(na2414_1), .EN(na252_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1701_1_i) );
// C_///AND/D      x135y34     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1702_4 ( .OUT(na1702_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1702_5 ( .OUT(na1702_2), .CLK(na2414_1), .EN(na253_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1702_2_i) );
// C_AND/D///      x138y33     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1703_1 ( .OUT(na1703_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1703_2 ( .OUT(na1703_1), .CLK(na2414_1), .EN(na253_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1703_1_i) );
// C_///AND/D      x132y47     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1704_4 ( .OUT(na1704_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1704_5 ( .OUT(na1704_2), .CLK(na2414_1), .EN(na253_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1704_2_i) );
// C_AND/D///      x137y48     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1705_1 ( .OUT(na1705_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1705_2 ( .OUT(na1705_1), .CLK(na2414_1), .EN(na253_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1705_1_i) );
// C_///AND/D      x135y70     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1706_4 ( .OUT(na1706_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1706_5 ( .OUT(na1706_2), .CLK(na2414_1), .EN(na253_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1706_2_i) );
// C_///AND/D      x133y63     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1707_4 ( .OUT(na1707_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2406_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1707_5 ( .OUT(na1707_2), .CLK(na2414_1), .EN(na253_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1707_2_i) );
// C_///AND/D      x132y70     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1708_4 ( .OUT(na1708_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1708_5 ( .OUT(na1708_2), .CLK(na2414_1), .EN(na253_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1708_2_i) );
// C_AND/D///      x135y70     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1709_1 ( .OUT(na1709_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1709_2 ( .OUT(na1709_1), .CLK(na2414_1), .EN(na253_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1709_1_i) );
// C_///AND/D      x138y82     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1710_4 ( .OUT(na1710_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1710_5 ( .OUT(na1710_2), .CLK(na2414_1), .EN(na253_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1710_2_i) );
// C_AND/D///      x152y81     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1711_1 ( .OUT(na1711_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1711_2 ( .OUT(na1711_1), .CLK(na2414_1), .EN(na253_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1711_1_i) );
// C_///AND/D      x155y32     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1712_4 ( .OUT(na1712_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1712_5 ( .OUT(na1712_2), .CLK(na2414_1), .EN(na248_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1712_2_i) );
// C_AND/D///      x140y35     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1713_1 ( .OUT(na1713_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1713_2 ( .OUT(na1713_1), .CLK(na2414_1), .EN(na248_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1713_1_i) );
// C_AND/D///      x126y43     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1714_1 ( .OUT(na1714_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2403_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1714_2 ( .OUT(na1714_1), .CLK(na2414_1), .EN(na248_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1714_1_i) );
// C_AND/D///      x138y47     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1715_1 ( .OUT(na1715_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1715_2 ( .OUT(na1715_1), .CLK(na2414_1), .EN(na248_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1715_1_i) );
// C_///AND/D      x137y72     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1716_4 ( .OUT(na1716_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1716_5 ( .OUT(na1716_2), .CLK(na2414_1), .EN(na248_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1716_2_i) );
// C_AND/D///      x138y63     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1717_1 ( .OUT(na1717_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1717_2 ( .OUT(na1717_1), .CLK(na2414_1), .EN(na248_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1717_1_i) );
// C_///AND/D      x131y75     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1718_4 ( .OUT(na1718_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1718_5 ( .OUT(na1718_2), .CLK(na2414_1), .EN(na248_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1718_2_i) );
// C_AND/D///      x134y72     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1719_1 ( .OUT(na1719_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1719_2 ( .OUT(na1719_1), .CLK(na2414_1), .EN(na248_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1719_1_i) );
// C_///AND/D      x138y76     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1720_4 ( .OUT(na1720_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1720_5 ( .OUT(na1720_2), .CLK(na2414_1), .EN(na248_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1720_2_i) );
// C_///AND/D      x142y83     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1721_4 ( .OUT(na1721_2_i), .IN1(1'b1), .IN2(na2410_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1721_5 ( .OUT(na1721_2), .CLK(na2414_1), .EN(na248_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1721_2_i) );
// C_///AND/D      x156y36     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1722_4 ( .OUT(na1722_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1722_5 ( .OUT(na1722_2), .CLK(na2414_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1722_2_i) );
// C_AND/D///      x140y36     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1723_1 ( .OUT(na1723_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1723_2 ( .OUT(na1723_1), .CLK(na2414_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1723_1_i) );
// C_///AND/D      x146y48     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1724_4 ( .OUT(na1724_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1724_5 ( .OUT(na1724_2), .CLK(na2414_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1724_2_i) );
// C_AND/D///      x145y45     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1725_1 ( .OUT(na1725_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1725_2 ( .OUT(na1725_1), .CLK(na2414_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1725_1_i) );
// C_///AND/D      x154y57     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1726_4 ( .OUT(na1726_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1726_5 ( .OUT(na1726_2), .CLK(na2414_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1726_2_i) );
// C_AND/D///      x153y63     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1727_1 ( .OUT(na1727_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1727_2 ( .OUT(na1727_1), .CLK(na2414_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1727_1_i) );
// C_AND/D///      x150y67     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1728_1 ( .OUT(na1728_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2407_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1728_2 ( .OUT(na1728_1), .CLK(na2414_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1728_1_i) );
// C_AND/D///      x156y69     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1729_1 ( .OUT(na1729_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1729_2 ( .OUT(na1729_1), .CLK(na2414_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1729_1_i) );
// C_///AND/D      x156y79     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1730_4 ( .OUT(na1730_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1730_5 ( .OUT(na1730_2), .CLK(na2414_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1730_2_i) );
// C_AND/D///      x140y81     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1731_1 ( .OUT(na1731_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1731_2 ( .OUT(na1731_1), .CLK(na2414_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1731_1_i) );
// C_///AND/D      x151y40     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1732_4 ( .OUT(na1732_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1732_5 ( .OUT(na1732_2), .CLK(na2414_1), .EN(na257_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1732_2_i) );
// C_AND/D///      x143y38     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1733_1 ( .OUT(na1733_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1733_2 ( .OUT(na1733_1), .CLK(na2414_1), .EN(na257_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1733_1_i) );
// C_///AND/D      x147y46     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1734_4 ( .OUT(na1734_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1734_5 ( .OUT(na1734_2), .CLK(na2414_1), .EN(na257_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1734_2_i) );
// C_///AND/D      x132y46     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1735_4 ( .OUT(na1735_2_i), .IN1(1'b1), .IN2(na2404_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1735_5 ( .OUT(na1735_2), .CLK(na2414_1), .EN(na257_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1735_2_i) );
// C_///AND/D      x151y54     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1736_4 ( .OUT(na1736_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1736_5 ( .OUT(na1736_2), .CLK(na2414_1), .EN(na257_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1736_2_i) );
// C_AND/D///      x151y59     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1737_1 ( .OUT(na1737_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1737_2 ( .OUT(na1737_1), .CLK(na2414_1), .EN(na257_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1737_1_i) );
// C_///AND/D      x144y67     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1738_4 ( .OUT(na1738_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1738_5 ( .OUT(na1738_2), .CLK(na2414_1), .EN(na257_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1738_2_i) );
// C_AND/D///      x149y66     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1739_1 ( .OUT(na1739_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1739_2 ( .OUT(na1739_1), .CLK(na2414_1), .EN(na257_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1739_1_i) );
// C_///AND/D      x153y69     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1740_4 ( .OUT(na1740_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1740_5 ( .OUT(na1740_2), .CLK(na2414_1), .EN(na257_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1740_2_i) );
// C_AND/D///      x138y79     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1741_1 ( .OUT(na1741_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1741_2 ( .OUT(na1741_1), .CLK(na2414_1), .EN(na257_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1741_1_i) );
// C_AND/D///      x154y35     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1742_1 ( .OUT(na1742_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2401_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1742_2 ( .OUT(na1742_1), .CLK(na2414_1), .EN(na258_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1742_1_i) );
// C_AND/D///      x144y39     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1743_1 ( .OUT(na1743_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1743_2 ( .OUT(na1743_1), .CLK(na2414_1), .EN(na258_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1743_1_i) );
// C_///AND/D      x144y47     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1744_4 ( .OUT(na1744_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1744_5 ( .OUT(na1744_2), .CLK(na2414_1), .EN(na258_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1744_2_i) );
// C_AND/D///      x141y41     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1745_1 ( .OUT(na1745_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1745_2 ( .OUT(na1745_1), .CLK(na2414_1), .EN(na258_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1745_1_i) );
// C_///AND/D      x152y53     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1746_4 ( .OUT(na1746_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1746_5 ( .OUT(na1746_2), .CLK(na2414_1), .EN(na258_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1746_2_i) );
// C_AND/D///      x148y60     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1747_1 ( .OUT(na1747_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1747_2 ( .OUT(na1747_1), .CLK(na2414_1), .EN(na258_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1747_1_i) );
// C_///AND/D      x147y70     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1748_4 ( .OUT(na1748_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1748_5 ( .OUT(na1748_2), .CLK(na2414_1), .EN(na258_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1748_2_i) );
// C_///AND/D      x156y65     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1749_4 ( .OUT(na1749_2_i), .IN1(na2408_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1749_5 ( .OUT(na1749_2), .CLK(na2414_1), .EN(na258_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1749_2_i) );
// C_///AND/D      x156y72     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1750_4 ( .OUT(na1750_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1750_5 ( .OUT(na1750_2), .CLK(na2414_1), .EN(na258_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1750_2_i) );
// C_AND/D///      x139y80     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1751_1 ( .OUT(na1751_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1751_2 ( .OUT(na1751_1), .CLK(na2414_1), .EN(na258_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1751_1_i) );
// C_///AND/D      x150y42     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1752_4 ( .OUT(na1752_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1752_5 ( .OUT(na1752_2), .CLK(na2414_1), .EN(na259_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1752_2_i) );
// C_AND/D///      x140y40     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1753_1 ( .OUT(na1753_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1753_2 ( .OUT(na1753_1), .CLK(na2414_1), .EN(na259_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1753_1_i) );
// C_///AND/D      x146y46     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1754_4 ( .OUT(na1754_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1754_5 ( .OUT(na1754_2), .CLK(na2414_1), .EN(na259_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1754_2_i) );
// C_AND/D///      x143y42     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1755_1 ( .OUT(na1755_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1755_2 ( .OUT(na1755_1), .CLK(na2414_1), .EN(na259_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1755_1_i) );
// C_AND/D///      x154y46     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1756_1 ( .OUT(na1756_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2405_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1756_2 ( .OUT(na1756_1), .CLK(na2414_1), .EN(na259_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1756_1_i) );
// C_AND/D///      x150y59     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1757_1 ( .OUT(na1757_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1757_2 ( .OUT(na1757_1), .CLK(na2414_1), .EN(na259_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1757_1_i) );
// C_///AND/D      x143y69     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1758_4 ( .OUT(na1758_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1758_5 ( .OUT(na1758_2), .CLK(na2414_1), .EN(na259_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1758_2_i) );
// C_AND/D///      x152y68     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1759_1 ( .OUT(na1759_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1759_2 ( .OUT(na1759_1), .CLK(na2414_1), .EN(na259_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1759_1_i) );
// C_///AND/D      x156y71     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1760_4 ( .OUT(na1760_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1760_5 ( .OUT(na1760_2), .CLK(na2414_1), .EN(na259_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1760_2_i) );
// C_AND/D///      x141y79     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1761_1 ( .OUT(na1761_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1761_2 ( .OUT(na1761_1), .CLK(na2414_1), .EN(na259_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1761_1_i) );
// C_///AND/D      x153y39     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1762_4 ( .OUT(na1762_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1762_5 ( .OUT(na1762_2), .CLK(na2414_1), .EN(na260_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1762_2_i) );
// C_///AND/D      x137y39     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1763_4 ( .OUT(na1763_2_i), .IN1(na2402_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1763_5 ( .OUT(na1763_2), .CLK(na2414_1), .EN(na260_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1763_2_i) );
// C_///AND/D      x142y40     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1764_4 ( .OUT(na1764_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1764_5 ( .OUT(na1764_2), .CLK(na2414_1), .EN(na260_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1764_2_i) );
// C_AND/D///      x141y46     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1765_1 ( .OUT(na1765_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1765_2 ( .OUT(na1765_1), .CLK(na2414_1), .EN(na260_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1765_1_i) );
// C_///AND/D      x153y55     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1766_4 ( .OUT(na1766_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1766_5 ( .OUT(na1766_2), .CLK(na2414_1), .EN(na260_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1766_2_i) );
// C_AND/D///      x151y63     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1767_1 ( .OUT(na1767_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1767_2 ( .OUT(na1767_1), .CLK(na2414_1), .EN(na260_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1767_1_i) );
// C_///AND/D      x148y65     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1768_4 ( .OUT(na1768_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1768_5 ( .OUT(na1768_2), .CLK(na2414_1), .EN(na260_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1768_2_i) );
// C_AND/D///      x153y65     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1769_1 ( .OUT(na1769_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1769_2 ( .OUT(na1769_1), .CLK(na2414_1), .EN(na260_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1769_1_i) );
// C_AND/D///      x153y79     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1770_1 ( .OUT(na1770_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2409_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1770_2 ( .OUT(na1770_1), .CLK(na2414_1), .EN(na260_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1770_1_i) );
// C_AND/D///      x139y73     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1771_1 ( .OUT(na1771_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1771_2 ( .OUT(na1771_1), .CLK(na2414_1), .EN(na260_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1771_1_i) );
// C_///AND/D      x155y40     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1772_4 ( .OUT(na1772_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1772_5 ( .OUT(na1772_2), .CLK(na2414_1), .EN(na261_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1772_2_i) );
// C_AND/D///      x137y40     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1773_1 ( .OUT(na1773_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1773_2 ( .OUT(na1773_1), .CLK(na2414_1), .EN(na261_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1773_1_i) );
// C_///AND/D      x144y41     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1774_4 ( .OUT(na1774_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1774_5 ( .OUT(na1774_2), .CLK(na2414_1), .EN(na261_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1774_2_i) );
// C_AND/D///      x143y45     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1775_1 ( .OUT(na1775_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1775_2 ( .OUT(na1775_1), .CLK(na2414_1), .EN(na261_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1775_1_i) );
// C_///AND/D      x155y56     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1776_4 ( .OUT(na1776_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1776_5 ( .OUT(na1776_2), .CLK(na2414_1), .EN(na261_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1776_2_i) );
// C_///AND/D      x147y66     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1777_4 ( .OUT(na1777_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2406_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1777_5 ( .OUT(na1777_2), .CLK(na2414_1), .EN(na261_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1777_2_i) );
// C_///AND/D      x152y66     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1778_4 ( .OUT(na1778_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1778_5 ( .OUT(na1778_2), .CLK(na2414_1), .EN(na261_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1778_2_i) );
// C_AND/D///      x153y68     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1779_1 ( .OUT(na1779_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1779_2 ( .OUT(na1779_1), .CLK(na2414_1), .EN(na261_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1779_1_i) );
// C_///AND/D      x155y80     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1780_4 ( .OUT(na1780_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1780_5 ( .OUT(na1780_2), .CLK(na2414_1), .EN(na261_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1780_2_i) );
// C_AND/D///      x141y74     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1781_1 ( .OUT(na1781_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1781_2 ( .OUT(na1781_1), .CLK(na2414_1), .EN(na261_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1781_1_i) );
// C_///AND/D      x156y43     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1782_4 ( .OUT(na1782_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1782_5 ( .OUT(na1782_2), .CLK(na2414_1), .EN(na262_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1782_2_i) );
// C_AND/D///      x140y39     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1783_1 ( .OUT(na1783_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1783_2 ( .OUT(na1783_1), .CLK(na2414_1), .EN(na262_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1783_1_i) );
// C_AND/D///      x153y38     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1784_1 ( .OUT(na1784_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2403_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1784_2 ( .OUT(na1784_1), .CLK(na2414_1), .EN(na262_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1784_1_i) );
// C_AND/D///      x140y44     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1785_1 ( .OUT(na1785_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1785_2 ( .OUT(na1785_1), .CLK(na2414_1), .EN(na262_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1785_1_i) );
// C_///AND/D      x156y57     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1786_4 ( .OUT(na1786_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1786_5 ( .OUT(na1786_2), .CLK(na2414_1), .EN(na262_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1786_2_i) );
// C_AND/D///      x152y63     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1787_1 ( .OUT(na1787_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1787_2 ( .OUT(na1787_1), .CLK(na2414_1), .EN(na262_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1787_1_i) );
// C_///AND/D      x149y67     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1788_4 ( .OUT(na1788_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1788_5 ( .OUT(na1788_2), .CLK(na2414_1), .EN(na262_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1788_2_i) );
// C_AND/D///      x154y67     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1789_1 ( .OUT(na1789_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1789_2 ( .OUT(na1789_1), .CLK(na2414_1), .EN(na262_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1789_1_i) );
// C_///AND/D      x148y83     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1790_4 ( .OUT(na1790_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1790_5 ( .OUT(na1790_2), .CLK(na2414_1), .EN(na262_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1790_2_i) );
// C_///AND/D      x136y83     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1791_4 ( .OUT(na1791_2_i), .IN1(1'b1), .IN2(na2410_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1791_5 ( .OUT(na1791_2), .CLK(na2414_1), .EN(na262_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1791_2_i) );
// C_///AND/D      x156y44     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1792_4 ( .OUT(na1792_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1792_5 ( .OUT(na1792_2), .CLK(na2414_1), .EN(na263_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1792_2_i) );
// C_AND/D///      x140y38     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1793_1 ( .OUT(na1793_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1793_2 ( .OUT(na1793_1), .CLK(na2414_1), .EN(na263_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1793_1_i) );
// C_///AND/D      x147y43     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1794_4 ( .OUT(na1794_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1794_5 ( .OUT(na1794_2), .CLK(na2414_1), .EN(na263_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1794_2_i) );
// C_AND/D///      x146y45     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1795_1 ( .OUT(na1795_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1795_2 ( .OUT(na1795_1), .CLK(na2414_1), .EN(na263_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1795_1_i) );
// C_///AND/D      x152y58     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1796_4 ( .OUT(na1796_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1796_5 ( .OUT(na1796_2), .CLK(na2414_1), .EN(na263_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1796_2_i) );
// C_AND/D///      x152y64     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1797_1 ( .OUT(na1797_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1797_2 ( .OUT(na1797_1), .CLK(na2414_1), .EN(na263_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1797_1_i) );
// C_AND/D///      x149y64     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1798_1 ( .OUT(na1798_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2407_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1798_2 ( .OUT(na1798_1), .CLK(na2414_1), .EN(na263_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1798_1_i) );
// C_AND/D///      x154y68     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1799_1 ( .OUT(na1799_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1799_2 ( .OUT(na1799_1), .CLK(na2414_1), .EN(na263_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1799_1_i) );
// C_///AND/D      x152y82     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1800_4 ( .OUT(na1800_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1800_5 ( .OUT(na1800_2), .CLK(na2414_1), .EN(na263_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1800_2_i) );
// C_AND/D///      x140y76     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1801_1 ( .OUT(na1801_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1801_2 ( .OUT(na1801_1), .CLK(na2414_1), .EN(na263_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1801_1_i) );
// C_///AND/D      x152y35     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1802_4 ( .OUT(na1802_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1802_5 ( .OUT(na1802_2), .CLK(na2414_1), .EN(na264_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1802_2_i) );
// C_AND/D///      x140y33     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1803_1 ( .OUT(na1803_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1803_2 ( .OUT(na1803_1), .CLK(na2414_1), .EN(na264_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1803_1_i) );
// C_///AND/D      x146y44     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1804_4 ( .OUT(na1804_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1804_5 ( .OUT(na1804_2), .CLK(na2414_1), .EN(na264_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1804_2_i) );
// C_///AND/D      x132y43     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1805_4 ( .OUT(na1805_2_i), .IN1(1'b1), .IN2(na2404_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1805_5 ( .OUT(na1805_2), .CLK(na2414_1), .EN(na264_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1805_2_i) );
// C_///AND/D      x151y60     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1806_4 ( .OUT(na1806_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1806_5 ( .OUT(na1806_2), .CLK(na2414_1), .EN(na264_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1806_2_i) );
// C_AND/D///      x150y62     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1807_1 ( .OUT(na1807_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1807_2 ( .OUT(na1807_1), .CLK(na2414_1), .EN(na264_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1807_1_i) );
// C_///AND/D      x148y68     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1808_4 ( .OUT(na1808_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1808_5 ( .OUT(na1808_2), .CLK(na2414_1), .EN(na264_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1808_2_i) );
// C_AND/D///      x151y69     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1809_1 ( .OUT(na1809_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1809_2 ( .OUT(na1809_1), .CLK(na2414_1), .EN(na264_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1809_1_i) );
// C_///AND/D      x153y74     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1810_4 ( .OUT(na1810_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1810_5 ( .OUT(na1810_2), .CLK(na2414_1), .EN(na264_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1810_2_i) );
// C_AND/D///      x137y75     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1811_1 ( .OUT(na1811_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1811_2 ( .OUT(na1811_1), .CLK(na2414_1), .EN(na264_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1811_1_i) );
// C_AND/D///      x153y35     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1812_1 ( .OUT(na1812_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2401_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1812_2 ( .OUT(na1812_1), .CLK(na2414_1), .EN(na255_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1812_1_i) );
// C_AND/D///      x141y39     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1813_1 ( .OUT(na1813_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1813_2 ( .OUT(na1813_1), .CLK(na2414_1), .EN(na255_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1813_1_i) );
// C_///AND/D      x147y49     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1814_4 ( .OUT(na1814_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1814_5 ( .OUT(na1814_2), .CLK(na2414_1), .EN(na255_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1814_2_i) );
// C_AND/D///      x142y43     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1815_1 ( .OUT(na1815_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1815_2 ( .OUT(na1815_1), .CLK(na2414_1), .EN(na255_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1815_1_i) );
// C_///AND/D      x153y53     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1816_4 ( .OUT(na1816_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1816_5 ( .OUT(na1816_2), .CLK(na2414_1), .EN(na255_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1816_2_i) );
// C_AND/D///      x149y60     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1817_1 ( .OUT(na1817_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1817_2 ( .OUT(na1817_1), .CLK(na2414_1), .EN(na255_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1817_1_i) );
// C_///AND/D      x146y70     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1818_4 ( .OUT(na1818_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1818_5 ( .OUT(na1818_2), .CLK(na2414_1), .EN(na255_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1818_2_i) );
// C_///AND/D      x155y65     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1819_4 ( .OUT(na1819_2_i), .IN1(na2408_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1819_5 ( .OUT(na1819_2), .CLK(na2414_1), .EN(na255_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1819_2_i) );
// C_///AND/D      x155y74     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1820_4 ( .OUT(na1820_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1820_5 ( .OUT(na1820_2), .CLK(na2414_1), .EN(na255_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1820_2_i) );
// C_AND/D///      x140y80     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1821_1 ( .OUT(na1821_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1821_2 ( .OUT(na1821_1), .CLK(na2414_1), .EN(na255_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1821_1_i) );
// C_///AND/D      x149y37     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1822_4 ( .OUT(na1822_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1822_5 ( .OUT(na1822_2), .CLK(na2414_1), .EN(na266_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1822_2_i) );
// C_AND/D///      x141y33     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1823_1 ( .OUT(na1823_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1823_2 ( .OUT(na1823_1), .CLK(na2414_1), .EN(na266_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1823_1_i) );
// C_///AND/D      x149y46     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1824_4 ( .OUT(na1824_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1824_5 ( .OUT(na1824_2), .CLK(na2414_1), .EN(na266_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1824_2_i) );
// C_AND/D///      x145y41     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1825_1 ( .OUT(na1825_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1825_2 ( .OUT(na1825_1), .CLK(na2414_1), .EN(na266_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1825_1_i) );
// C_AND/D///      x156y48     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1826_1 ( .OUT(na1826_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2405_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1826_2 ( .OUT(na1826_1), .CLK(na2414_1), .EN(na266_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1826_1_i) );
// C_AND/D///      x151y62     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1827_1 ( .OUT(na1827_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1827_2 ( .OUT(na1827_1), .CLK(na2414_1), .EN(na266_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1827_1_i) );
// C_///AND/D      x151y72     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1828_4 ( .OUT(na1828_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1828_5 ( .OUT(na1828_2), .CLK(na2414_1), .EN(na266_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1828_2_i) );
// C_AND/D///      x152y67     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1829_1 ( .OUT(na1829_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1829_2 ( .OUT(na1829_1), .CLK(na2414_1), .EN(na266_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1829_1_i) );
// C_///AND/D      x156y74     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1830_4 ( .OUT(na1830_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1830_5 ( .OUT(na1830_2), .CLK(na2414_1), .EN(na266_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1830_2_i) );
// C_AND/D///      x140y77     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1831_1 ( .OUT(na1831_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1831_2 ( .OUT(na1831_1), .CLK(na2414_1), .EN(na266_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1831_1_i) );
// C_///AND/D      x151y38     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1832_4 ( .OUT(na1832_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1832_5 ( .OUT(na1832_2), .CLK(na2414_1), .EN(na267_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1832_2_i) );
// C_///AND/D      x137y42     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1833_4 ( .OUT(na1833_2_i), .IN1(na2402_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1833_5 ( .OUT(na1833_2), .CLK(na2414_1), .EN(na267_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1833_2_i) );
// C_///AND/D      x151y45     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1834_4 ( .OUT(na1834_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1834_5 ( .OUT(na1834_2), .CLK(na2414_1), .EN(na267_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1834_2_i) );
// C_AND/D///      x145y44     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1835_1 ( .OUT(na1835_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1835_2 ( .OUT(na1835_1), .CLK(na2414_1), .EN(na267_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1835_1_i) );
// C_///AND/D      x152y59     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1836_4 ( .OUT(na1836_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1836_5 ( .OUT(na1836_2), .CLK(na2414_1), .EN(na267_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1836_2_i) );
// C_AND/D///      x151y61     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1837_1 ( .OUT(na1837_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1837_2 ( .OUT(na1837_1), .CLK(na2414_1), .EN(na267_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1837_1_i) );
// C_///AND/D      x149y73     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1838_4 ( .OUT(na1838_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1838_5 ( .OUT(na1838_2), .CLK(na2414_1), .EN(na267_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1838_2_i) );
// C_AND/D///      x154y72     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1839_1 ( .OUT(na1839_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1839_2 ( .OUT(na1839_1), .CLK(na2414_1), .EN(na267_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1839_1_i) );
// C_AND/D///      x154y79     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1840_1 ( .OUT(na1840_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2409_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1840_2 ( .OUT(na1840_1), .CLK(na2414_1), .EN(na267_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1840_1_i) );
// C_AND/D///      x140y78     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1841_1 ( .OUT(na1841_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1841_2 ( .OUT(na1841_1), .CLK(na2414_1), .EN(na267_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1841_1_i) );
// C_///AND/D      x155y35     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1842_4 ( .OUT(na1842_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1842_5 ( .OUT(na1842_2), .CLK(na2414_1), .EN(na268_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1842_2_i) );
// C_AND/D///      x141y37     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1843_1 ( .OUT(na1843_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1843_2 ( .OUT(na1843_1), .CLK(na2414_1), .EN(na268_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1843_1_i) );
// C_///AND/D      x149y49     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1844_4 ( .OUT(na1844_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1844_5 ( .OUT(na1844_2), .CLK(na2414_1), .EN(na268_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1844_2_i) );
// C_AND/D///      x148y48     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1845_1 ( .OUT(na1845_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1845_2 ( .OUT(na1845_1), .CLK(na2414_1), .EN(na268_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1845_1_i) );
// C_///AND/D      x153y60     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1846_4 ( .OUT(na1846_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1846_5 ( .OUT(na1846_2), .CLK(na2414_1), .EN(na268_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1846_2_i) );
// C_///AND/D      x156y64     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1847_4 ( .OUT(na1847_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2406_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1847_5 ( .OUT(na1847_2), .CLK(na2414_1), .EN(na268_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1847_2_i) );
// C_///AND/D      x147y72     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1848_4 ( .OUT(na1848_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1848_5 ( .OUT(na1848_2), .CLK(na2414_1), .EN(na268_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1848_2_i) );
// C_AND/D///      x153y72     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1849_1 ( .OUT(na1849_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1849_2 ( .OUT(na1849_1), .CLK(na2414_1), .EN(na268_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1849_1_i) );
// C_///AND/D      x151y82     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1850_4 ( .OUT(na1850_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1850_5 ( .OUT(na1850_2), .CLK(na2414_1), .EN(na268_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1850_2_i) );
// C_AND/D///      x141y84     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1851_1 ( .OUT(na1851_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1851_2 ( .OUT(na1851_1), .CLK(na2414_1), .EN(na268_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1851_1_i) );
// C_///AND/D      x155y38     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1852_4 ( .OUT(na1852_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1852_5 ( .OUT(na1852_2), .CLK(na2414_1), .EN(na269_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1852_2_i) );
// C_AND/D///      x139y38     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1853_1 ( .OUT(na1853_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1853_2 ( .OUT(na1853_1), .CLK(na2414_1), .EN(na269_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1853_1_i) );
// C_AND/D///      x153y40     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1854_1 ( .OUT(na1854_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2403_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1854_2 ( .OUT(na1854_1), .CLK(na2414_1), .EN(na269_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1854_1_i) );
// C_AND/D///      x146y47     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1855_1 ( .OUT(na1855_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1855_2 ( .OUT(na1855_1), .CLK(na2414_1), .EN(na269_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1855_1_i) );
// C_///AND/D      x155y59     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1856_4 ( .OUT(na1856_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1856_5 ( .OUT(na1856_2), .CLK(na2414_1), .EN(na269_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1856_2_i) );
// C_AND/D///      x154y63     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1857_1 ( .OUT(na1857_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1857_2 ( .OUT(na1857_1), .CLK(na2414_1), .EN(na269_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1857_1_i) );
// C_///AND/D      x149y69     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1858_4 ( .OUT(na1858_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1858_5 ( .OUT(na1858_2), .CLK(na2414_1), .EN(na269_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1858_2_i) );
// C_AND/D///      x153y71     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1859_1 ( .OUT(na1859_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1859_2 ( .OUT(na1859_1), .CLK(na2414_1), .EN(na269_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1859_1_i) );
// C_///AND/D      x153y81     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1860_4 ( .OUT(na1860_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1860_5 ( .OUT(na1860_2), .CLK(na2414_1), .EN(na269_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1860_2_i) );
// C_///AND/D      x139y83     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1861_4 ( .OUT(na1861_2_i), .IN1(1'b1), .IN2(na2410_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1861_5 ( .OUT(na1861_2), .CLK(na2414_1), .EN(na269_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1861_2_i) );
// C_///AND/D      x154y37     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1862_4 ( .OUT(na1862_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1862_5 ( .OUT(na1862_2), .CLK(na2414_1), .EN(na270_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1862_2_i) );
// C_AND/D///      x140y37     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1863_1 ( .OUT(na1863_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1863_2 ( .OUT(na1863_1), .CLK(na2414_1), .EN(na270_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1863_1_i) );
// C_///AND/D      x154y49     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1864_4 ( .OUT(na1864_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1864_5 ( .OUT(na1864_2), .CLK(na2414_1), .EN(na270_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1864_2_i) );
// C_AND/D///      x147y48     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1865_1 ( .OUT(na1865_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1865_2 ( .OUT(na1865_1), .CLK(na2414_1), .EN(na270_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1865_1_i) );
// C_///AND/D      x156y60     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1866_4 ( .OUT(na1866_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1866_5 ( .OUT(na1866_2), .CLK(na2414_1), .EN(na270_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1866_2_i) );
// C_AND/D///      x151y64     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1867_1 ( .OUT(na1867_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1867_2 ( .OUT(na1867_1), .CLK(na2414_1), .EN(na270_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1867_1_i) );
// C_AND/D///      x150y68     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1868_1 ( .OUT(na1868_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2407_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1868_2 ( .OUT(na1868_1), .CLK(na2414_1), .EN(na270_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1868_1_i) );
// C_AND/D///      x154y70     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1869_1 ( .OUT(na1869_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1869_2 ( .OUT(na1869_1), .CLK(na2414_1), .EN(na270_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1869_1_i) );
// C_///AND/D      x156y82     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1870_4 ( .OUT(na1870_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1870_5 ( .OUT(na1870_2), .CLK(na2414_1), .EN(na270_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1870_2_i) );
// C_AND/D///      x140y82     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1871_1 ( .OUT(na1871_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1871_2 ( .OUT(na1871_1), .CLK(na2414_1), .EN(na270_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1871_1_i) );
// C_///AND/D      x148y38     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1872_4 ( .OUT(na1872_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2401_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1872_5 ( .OUT(na1872_2), .CLK(na2414_1), .EN(na265_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1872_2_i) );
// C_AND/D///      x140y34     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1873_1 ( .OUT(na1873_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2402_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1873_2 ( .OUT(na1873_1), .CLK(na2414_1), .EN(na265_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1873_1_i) );
// C_///AND/D      x148y47     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1874_4 ( .OUT(na1874_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2403_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1874_5 ( .OUT(na1874_2), .CLK(na2414_1), .EN(na265_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1874_2_i) );
// C_///AND/D      x138y48     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1875_4 ( .OUT(na1875_2_i), .IN1(1'b1), .IN2(na2404_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1875_5 ( .OUT(na1875_2), .CLK(na2414_1), .EN(na265_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1875_2_i) );
// C_///AND/D      x155y63     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1876_4 ( .OUT(na1876_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2405_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1876_5 ( .OUT(na1876_2), .CLK(na2414_1), .EN(na265_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1876_2_i) );
// C_AND/D///      x150y63     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1877_1 ( .OUT(na1877_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2406_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1877_2 ( .OUT(na1877_1), .CLK(na2414_1), .EN(na265_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1877_1_i) );
// C_///AND/D      x154y71     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1878_4 ( .OUT(na1878_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1878_5 ( .OUT(na1878_2), .CLK(na2414_1), .EN(na265_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1878_2_i) );
// C_AND/D///      x149y70     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1879_1 ( .OUT(na1879_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2408_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1879_2 ( .OUT(na1879_1), .CLK(na2414_1), .EN(na265_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1879_1_i) );
// C_///AND/D      x155y75     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1880_4 ( .OUT(na1880_2_i), .IN1(na2409_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1880_5 ( .OUT(na1880_2), .CLK(na2414_1), .EN(na265_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1880_2_i) );
// C_AND/D///      x139y78     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1881_1 ( .OUT(na1881_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1881_2 ( .OUT(na1881_1), .CLK(na2414_1), .EN(na265_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1881_1_i) );
// C_MX4b////      x146y36     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1882_1 ( .OUT(na1882_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na362_2), .IN6(na422_1), .IN7(na412_2),
                      .IN8(na352_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x146y37     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1883_1 ( .OUT(na1883_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na382_2), .IN6(na392_2), .IN7(na342_1),
                      .IN8(na282_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x149y38     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1884_1 ( .OUT(na1884_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na332_2), .IN6(na322_2), .IN7(na372_1),
                      .IN8(na592_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x145y37     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1885_1 ( .OUT(na1885_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na312_1), .IN6(na302_2), .IN7(na292_2),
                      .IN8(na432_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x145y38     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1886_1 ( .OUT(na1886_1), .IN1(~na2384_1), .IN2(1'b1), .IN3(~na2385_1), .IN4(1'b1), .IN5(na1885_1), .IN6(na1884_1), .IN7(na1883_1),
                      .IN8(na1882_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x142y37     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1887_1 ( .OUT(na1887_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na423_1), .IN6(na363_1), .IN7(na353_2),
                      .IN8(na413_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x140y32     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1888_1 ( .OUT(na1888_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na283_1), .IN6(na343_1), .IN7(na393_1),
                      .IN8(na383_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x139y31     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1889_1 ( .OUT(na1889_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na373_1), .IN6(na593_1), .IN7(na333_1),
                      .IN8(na323_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x145y34     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1890_1 ( .OUT(na1890_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na313_1), .IN6(na303_1), .IN7(na293_1),
                      .IN8(na433_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x137y34     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1891_1 ( .OUT(na1891_1), .IN1(na2384_1), .IN2(1'b1), .IN3(~na2385_1), .IN4(1'b1), .IN5(na1889_1), .IN6(na1890_1), .IN7(na1887_1),
                      .IN8(na1888_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x147y38     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1892_1 ( .OUT(na1892_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na354_2), .IN6(na414_2), .IN7(na424_2),
                      .IN8(na364_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x145y39     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1893_1 ( .OUT(na1893_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na384_2), .IN6(na394_1), .IN7(na344_2),
                      .IN8(na284_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x144y42     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1894_1 ( .OUT(na1894_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na594_2), .IN6(na374_2), .IN7(na324_2),
                      .IN8(na334_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x148y39     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1895_1 ( .OUT(na1895_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na294_2), .IN6(na434_2), .IN7(na314_2),
                      .IN8(na304_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x143y44     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1896_1 ( .OUT(na1896_1), .IN1(~na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na1893_1), .IN6(na1892_1), .IN7(na1895_1),
                      .IN8(na1894_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x126y47     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1897_1 ( .OUT(na1897_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na365_1), .IN6(na425_1), .IN7(na415_1),
                      .IN8(na355_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x128y48     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1898_1 ( .OUT(na1898_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na345_2), .IN6(na285_1), .IN7(na385_1),
                      .IN8(na395_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x123y47     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1899_1 ( .OUT(na1899_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na335_1), .IN6(na325_1), .IN7(na375_2),
                      .IN8(na595_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x125y48     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1900_1 ( .OUT(na1900_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na315_1), .IN6(na305_1), .IN7(na295_2),
                      .IN8(na435_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x132y48     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1901_1 ( .OUT(na1901_1), .IN1(na2384_1), .IN2(1'b1), .IN3(~na2385_1), .IN4(1'b1), .IN5(na1899_1), .IN6(na1900_1), .IN7(na1897_1),
                      .IN8(na1898_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x147y47     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1902_1 ( .OUT(na1902_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na366_2), .IN6(na426_2), .IN7(na416_1),
                      .IN8(na356_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x149y48     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1903_1 ( .OUT(na1903_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na396_2), .IN6(na386_1), .IN7(na286_2),
                      .IN8(na346_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x150y47     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1904_1 ( .OUT(na1904_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na596_2), .IN6(na376_2), .IN7(na326_2),
                      .IN8(na336_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x152y48     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1905_1 ( .OUT(na1905_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na316_2), .IN6(na306_1), .IN7(na296_2),
                      .IN8(na436_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x147y50     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1906_1 ( .OUT(na1906_1), .IN1(na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na1902_1), .IN6(na1903_1), .IN7(na1904_1),
                      .IN8(na1905_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x144y51     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1907_1 ( .OUT(na1907_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na367_2), .IN6(na427_2), .IN7(na417_1),
                      .IN8(na357_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x142y50     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1908_1 ( .OUT(na1908_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na397_2), .IN6(na387_1), .IN7(na287_2),
                      .IN8(na347_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x145y51     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1909_1 ( .OUT(na1909_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na337_1), .IN6(na327_1), .IN7(na377_1),
                      .IN8(na597_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x147y54     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1910_1 ( .OUT(na1910_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na317_2), .IN6(na307_1), .IN7(na297_1),
                      .IN8(na437_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x141y54     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1911_1 ( .OUT(na1911_1), .IN1(na2384_1), .IN2(1'b1), .IN3(~na2385_1), .IN4(1'b1), .IN5(na1909_1), .IN6(na1910_1), .IN7(na1907_1),
                      .IN8(na1908_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x143y56     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1912_1 ( .OUT(na1912_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na418_2), .IN6(na358_2), .IN7(na368_2),
                      .IN8(na428_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x141y59     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1913_1 ( .OUT(na1913_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na388_2), .IN6(na398_2), .IN7(na348_2),
                      .IN8(na288_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x142y62     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1914_1 ( .OUT(na1914_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na338_2), .IN6(na328_1), .IN7(na378_1),
                      .IN8(na598_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x144y61     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1915_1 ( .OUT(na1915_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na318_2), .IN6(na308_2), .IN7(na298_1),
                      .IN8(na438_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x143y60     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1916_1 ( .OUT(na1916_1), .IN1(~na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na1913_1), .IN6(na1912_1), .IN7(na1915_1),
                      .IN8(na1914_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x141y67     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1917_1 ( .OUT(na1917_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na419_2), .IN6(na359_1), .IN7(na369_1),
                      .IN8(na429_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x141y66     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1918_1 ( .OUT(na1918_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na399_1), .IN6(na389_2), .IN7(na289_1),
                      .IN8(na349_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x142y65     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1919_1 ( .OUT(na1919_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na339_2), .IN6(na329_1), .IN7(na379_1),
                      .IN8(na599_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x140y68     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1920_1 ( .OUT(na1920_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na299_1), .IN6(na439_1), .IN7(na319_1),
                      .IN8(na309_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x137y68     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1921_1 ( .OUT(na1921_1), .IN1(na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na1917_1), .IN6(na1918_1), .IN7(na1919_1),
                      .IN8(na1920_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x147y73     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1922_1 ( .OUT(na1922_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na420_2), .IN6(na360_2), .IN7(na370_2),
                      .IN8(na430_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x145y74     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1923_1 ( .OUT(na1923_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na400_1), .IN6(na390_2), .IN7(na290_1),
                      .IN8(na350_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x142y71     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1924_1 ( .OUT(na1924_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na600_2), .IN6(na380_2), .IN7(na330_2),
                      .IN8(na340_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x148y76     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1925_1 ( .OUT(na1925_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na320_1), .IN6(na310_2), .IN7(na300_2),
                      .IN8(na440_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x143y72     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1926_1 ( .OUT(na1926_1), .IN1(na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na1922_1), .IN6(na1923_1), .IN7(na1924_1),
                      .IN8(na1925_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x131y79     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1927_1 ( .OUT(na1927_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na371_1), .IN6(na431_1), .IN7(na421_1),
                      .IN8(na361_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x131y76     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1928_1 ( .OUT(na1928_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na291_1), .IN6(na351_1), .IN7(na401_1),
                      .IN8(na391_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x128y81     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1929_1 ( .OUT(na1929_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na381_1), .IN6(na601_1), .IN7(na341_1),
                      .IN8(na331_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x132y76     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1930_1 ( .OUT(na1930_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na311_1), .IN6(na321_1), .IN7(na441_2),
                      .IN8(na301_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x132y74     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1931_1 ( .OUT(na1931_1), .IN1(na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na1927_1), .IN6(na1928_1), .IN7(na1929_1),
                      .IN8(na1930_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x145y33     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1932_1 ( .OUT(na1932_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na692_2), .IN6(na612_2), .IN7(na622_2),
                      .IN8(na632_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x147y36     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1933_1 ( .OUT(na1933_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na642_1), .IN6(na652_2), .IN7(na662_2),
                      .IN8(na672_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x148y35     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1934_1 ( .OUT(na1934_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na682_2), .IN6(na752_1), .IN7(na702_1),
                      .IN8(na712_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x150y36     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1935_1 ( .OUT(na1935_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na722_2), .IN6(na732_2), .IN7(na742_2),
                      .IN8(na602_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x145y40     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1936_1 ( .OUT(na1936_1), .IN1(na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na1932_1), .IN6(na1933_1), .IN7(na1934_1),
                      .IN8(na1935_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x143y32     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1937_1 ( .OUT(na1937_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na623_1), .IN6(na633_1), .IN7(na693_1),
                      .IN8(na613_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x145y31     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1938_1 ( .OUT(na1938_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na663_1), .IN6(na673_1), .IN7(na643_1),
                      .IN8(na653_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x154y32     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1939_1 ( .OUT(na1939_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na683_2), .IN6(na753_1), .IN7(na703_1),
                      .IN8(na713_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x150y33     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1940_1 ( .OUT(na1940_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na603_2), .IN6(na743_1), .IN7(na733_1),
                      .IN8(na723_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x152y34     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1941_1 ( .OUT(na1941_1), .IN1(~na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na1938_1), .IN6(na1937_1), .IN7(na1940_1),
                      .IN8(na1939_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x146y43     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1942_1 ( .OUT(na1942_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na694_1), .IN6(na614_1), .IN7(na624_2),
                      .IN8(na634_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x150y44     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1943_1 ( .OUT(na1943_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na674_2), .IN6(na664_1), .IN7(na654_2),
                      .IN8(na644_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x145y43     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1944_1 ( .OUT(na1944_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na714_2), .IN6(na704_2), .IN7(na754_2),
                      .IN8(na684_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x147y44     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1945_1 ( .OUT(na1945_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na744_2), .IN6(na604_2), .IN7(na724_1),
                      .IN8(na734_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x145y46     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1946_1 ( .OUT(na1946_1), .IN1(na2384_1), .IN2(1'b1), .IN3(~na2385_1), .IN4(1'b1), .IN5(na1944_1), .IN6(na1945_1), .IN7(na1942_1),
                      .IN8(na1943_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x131y49     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1947_1 ( .OUT(na1947_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na695_1), .IN6(na615_1), .IN7(na625_2),
                      .IN8(na635_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x131y52     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1948_1 ( .OUT(na1948_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na655_1), .IN6(na645_1), .IN7(na675_2),
                      .IN8(na665_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x132y51     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1949_1 ( .OUT(na1949_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na755_1), .IN6(na685_1), .IN7(na715_1),
                      .IN8(na705_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x134y54     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1950_1 ( .OUT(na1950_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na725_1), .IN6(na735_2), .IN7(na745_1),
                      .IN8(na605_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x133y52     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1951_1 ( .OUT(na1951_1), .IN1(na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na1947_1), .IN6(na1948_1), .IN7(na1949_1),
                      .IN8(na1950_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x153y42     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1952_1 ( .OUT(na1952_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na616_2), .IN6(na696_2), .IN7(na636_1),
                      .IN8(na626_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x151y41     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1953_1 ( .OUT(na1953_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na656_2), .IN6(na646_2), .IN7(na676_2),
                      .IN8(na666_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x154y44     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1954_1 ( .OUT(na1954_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na706_2), .IN6(na716_1), .IN7(na686_1),
                      .IN8(na756_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x152y43     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1955_1 ( .OUT(na1955_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na736_2), .IN6(na726_2), .IN7(na606_1),
                      .IN8(na746_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x151y44     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1956_1 ( .OUT(na1956_1), .IN1(~na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na1953_1), .IN6(na1952_1), .IN7(na1955_1),
                      .IN8(na1954_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x150y50     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1957_1 ( .OUT(na1957_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na697_2), .IN6(na617_2), .IN7(na627_1),
                      .IN8(na637_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x152y49     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1958_1 ( .OUT(na1958_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na647_2), .IN6(na657_1), .IN7(na667_1),
                      .IN8(na677_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x155y52     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1959_1 ( .OUT(na1959_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na687_1), .IN6(na757_2), .IN7(na707_1),
                      .IN8(na717_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x151y51     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1960_1 ( .OUT(na1960_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na737_1), .IN6(na727_2), .IN7(na607_1),
                      .IN8(na747_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x147y52     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1961_1 ( .OUT(na1961_1), .IN1(~na2384_1), .IN2(1'b1), .IN3(~na2385_1), .IN4(1'b1), .IN5(na1960_1), .IN6(na1959_1), .IN7(na1958_1),
                      .IN8(na1957_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x143y62     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1962_1 ( .OUT(na1962_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na698_2), .IN6(na618_2), .IN7(na628_1),
                      .IN8(na638_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x143y63     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1963_1 ( .OUT(na1963_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na658_1), .IN6(na648_2), .IN7(na678_2),
                      .IN8(na668_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x146y64     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1964_1 ( .OUT(na1964_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na688_2), .IN6(na758_2), .IN7(na708_1),
                      .IN8(na718_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x148y61     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1965_1 ( .OUT(na1965_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na728_2), .IN6(na738_1), .IN7(na748_2),
                      .IN8(na608_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x141y62     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1966_1 ( .OUT(na1966_1), .IN1(~na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na1963_1), .IN6(na1962_1), .IN7(na1965_1),
                      .IN8(na1964_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x146y72     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1967_1 ( .OUT(na1967_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na619_1), .IN6(na699_1), .IN7(na639_2),
                      .IN8(na629_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x146y69     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1968_1 ( .OUT(na1968_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na679_1), .IN6(na669_2), .IN7(na659_1),
                      .IN8(na649_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x145y70     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1969_1 ( .OUT(na1969_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na759_1), .IN6(na689_1), .IN7(na719_2),
                      .IN8(na709_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x141y69     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1970_1 ( .OUT(na1970_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na729_1), .IN6(na739_1), .IN7(na749_2),
                      .IN8(na609_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x145y68     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1971_1 ( .OUT(na1971_1), .IN1(~na2384_1), .IN2(1'b1), .IN3(~na2385_1), .IN4(1'b1), .IN5(na1970_1), .IN6(na1969_1), .IN7(na1968_1),
                      .IN8(na1967_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x151y76     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1972_1 ( .OUT(na1972_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na630_2), .IN6(na640_2), .IN7(na700_2),
                      .IN8(na620_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x151y77     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1973_1 ( .OUT(na1973_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na680_1), .IN6(na670_2), .IN7(na660_2),
                      .IN8(na650_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x148y78     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1974_1 ( .OUT(na1974_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na710_2), .IN6(na720_2), .IN7(na690_2),
                      .IN8(na760_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x150y79     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1975_1 ( .OUT(na1975_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na740_2), .IN6(na730_1), .IN7(na610_2),
                      .IN8(na750_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x149y78     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1976_1 ( .OUT(na1976_1), .IN1(~na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na1973_1), .IN6(na1972_1), .IN7(na1975_1),
                      .IN8(na1974_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x133y77     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1977_1 ( .OUT(na1977_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na621_1), .IN6(na701_1), .IN7(na641_1),
                      .IN8(na631_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x135y82     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1978_1 ( .OUT(na1978_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na651_1), .IN6(na661_2), .IN7(na671_1),
                      .IN8(na681_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x134y75     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1979_1 ( .OUT(na1979_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na691_2), .IN6(na761_1), .IN7(na711_1),
                      .IN8(na721_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x136y82     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1980_1 ( .OUT(na1980_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na731_1), .IN6(na741_2), .IN7(na751_1),
                      .IN8(na611_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x135y76     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1981_1 ( .OUT(na1981_1), .IN1(na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na1977_1), .IN6(na1978_1), .IN7(na1979_1),
                      .IN8(na1980_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x115y32     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1982_1 ( .OUT(na1982_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na772_2), .IN6(na852_2), .IN7(na792_2),
                      .IN8(na782_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x117y31     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1983_1 ( .OUT(na1983_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na832_2), .IN6(na822_2), .IN7(na812_1),
                      .IN8(na802_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x120y32     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1984_1 ( .OUT(na1984_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na912_2), .IN6(na842_2), .IN7(na872_2),
                      .IN8(na862_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x122y31     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1985_1 ( .OUT(na1985_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na762_2), .IN6(na902_2), .IN7(na892_1),
                      .IN8(na882_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x118y34     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1986_1 ( .OUT(na1986_1), .IN1(~na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na1983_1), .IN6(na1982_1), .IN7(na1985_1),
                      .IN8(na1984_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x118y37     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1987_1 ( .OUT(na1987_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na853_1), .IN6(na773_1), .IN7(na783_1),
                      .IN8(na793_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x120y38     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1988_1 ( .OUT(na1988_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na823_2), .IN6(na833_1), .IN7(na803_1),
                      .IN8(na813_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x123y45     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1989_1 ( .OUT(na1989_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na843_1), .IN6(na913_1), .IN7(na863_1),
                      .IN8(na873_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x125y42     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1990_1 ( .OUT(na1990_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na883_1), .IN6(na893_1), .IN7(na903_2),
                      .IN8(na763_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x125y44     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1991_1 ( .OUT(na1991_1), .IN1(na2384_1), .IN2(1'b1), .IN3(~na2385_1), .IN4(1'b1), .IN5(na1989_1), .IN6(na1990_1), .IN7(na1987_1),
                      .IN8(na1988_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x114y42     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1992_1 ( .OUT(na1992_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na784_2), .IN6(na794_2), .IN7(na854_2),
                      .IN8(na774_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x120y39     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1993_1 ( .OUT(na1993_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na824_2), .IN6(na834_1), .IN7(na804_1),
                      .IN8(na814_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x119y38     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1994_1 ( .OUT(na1994_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na864_2), .IN6(na874_2), .IN7(na844_2),
                      .IN8(na914_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x117y35     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1995_1 ( .OUT(na1995_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na894_2), .IN6(na884_1), .IN7(na764_2),
                      .IN8(na904_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x118y39     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1996_1 ( .OUT(na1996_1), .IN1(~na2384_1), .IN2(1'b1), .IN3(~na2385_1), .IN4(1'b1), .IN5(na1995_1), .IN6(na1994_1), .IN7(na1993_1),
                      .IN8(na1992_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x120y47     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1997_1 ( .OUT(na1997_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na785_2), .IN6(na795_1), .IN7(na855_1),
                      .IN8(na775_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x114y44     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1998_1 ( .OUT(na1998_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na805_1), .IN6(na815_2), .IN7(na825_1),
                      .IN8(na835_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x117y43     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1999_1 ( .OUT(na1999_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na865_1), .IN6(na875_1), .IN7(na845_2),
                      .IN8(na915_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x119y46     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2000_1 ( .OUT(na2000_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na885_1), .IN6(na895_2), .IN7(na905_1),
                      .IN8(na765_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x120y46     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2001_1 ( .OUT(na2001_1), .IN1(na2384_1), .IN2(1'b1), .IN3(~na2385_1), .IN4(1'b1), .IN5(na1999_1), .IN6(na2000_1), .IN7(na1997_1),
                      .IN8(na1998_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x116y51     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2002_1 ( .OUT(na2002_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na856_1), .IN6(na776_2), .IN7(na786_2),
                      .IN8(na796_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x114y46     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2003_1 ( .OUT(na2003_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na826_1), .IN6(na836_2), .IN7(na806_2),
                      .IN8(na816_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x111y49     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2004_1 ( .OUT(na2004_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na846_2), .IN6(na916_2), .IN7(na866_2),
                      .IN8(na876_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x115y52     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2005_1 ( .OUT(na2005_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na896_2), .IN6(na886_2), .IN7(na766_2),
                      .IN8(na906_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x116y50     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2006_1 ( .OUT(na2006_1), .IN1(na2384_1), .IN2(1'b1), .IN3(~na2385_1), .IN4(1'b1), .IN5(na2004_1), .IN6(na2005_1), .IN7(na2002_1),
                      .IN8(na2003_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x125y52     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2007_1 ( .OUT(na2007_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na787_1), .IN6(na797_1), .IN7(na857_1),
                      .IN8(na777_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x127y53     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2008_1 ( .OUT(na2008_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na827_1), .IN6(na837_2), .IN7(na807_2),
                      .IN8(na817_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x124y56     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2009_1 ( .OUT(na2009_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na917_2), .IN6(na847_1), .IN7(na877_1),
                      .IN8(na867_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x126y55     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2010_1 ( .OUT(na2010_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na897_1), .IN6(na887_1), .IN7(na767_1),
                      .IN8(na907_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x126y53     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2011_1 ( .OUT(na2011_1), .IN1(~na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na2008_1), .IN6(na2007_1), .IN7(na2010_1),
                      .IN8(na2009_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x127y67     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2012_1 ( .OUT(na2012_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na858_2), .IN6(na778_2), .IN7(na788_2),
                      .IN8(na798_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x127y64     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2013_1 ( .OUT(na2013_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na828_2), .IN6(na838_2), .IN7(na808_2),
                      .IN8(na818_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x130y67     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2014_1 ( .OUT(na2014_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na848_1), .IN6(na918_2), .IN7(na868_2),
                      .IN8(na878_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x130y66     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2015_1 ( .OUT(na2015_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na908_2), .IN6(na768_1), .IN7(na888_2),
                      .IN8(na898_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x127y66     80'h00_0018_00_0040_0C0F_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2016_1 ( .OUT(na2016_1), .IN1(na2012_1), .IN2(na2013_1), .IN3(na2014_1), .IN4(na2015_1), .IN5(na2384_1), .IN6(1'b1), .IN7(na2385_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x121y67     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2017_1 ( .OUT(na2017_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na789_1), .IN6(na799_1), .IN7(na859_2),
                      .IN8(na779_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x125y68     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2018_1 ( .OUT(na2018_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na819_1), .IN6(na809_1), .IN7(na839_1),
                      .IN8(na829_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x124y69     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2019_1 ( .OUT(na2019_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na849_1), .IN6(na919_1), .IN7(na869_1),
                      .IN8(na879_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x122y70     80'h00_0018_00_0040_0C0F_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2020_1 ( .OUT(na2020_1), .IN1(na899_1), .IN2(na889_2), .IN3(na769_1), .IN4(na909_1), .IN5(~na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x125y70     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2021_1 ( .OUT(na2021_1), .IN1(na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na2017_1), .IN6(na2018_1), .IN7(na2019_1),
                      .IN8(na2020_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x116y76     80'h00_0018_00_0040_0C0F_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2022_1 ( .OUT(na2022_1), .IN1(na780_2), .IN2(na860_2), .IN3(na800_2), .IN4(na790_1), .IN5(~na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x116y75     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2023_1 ( .OUT(na2023_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na830_2), .IN6(na840_1), .IN7(na810_2),
                      .IN8(na820_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x115y76     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2024_1 ( .OUT(na2024_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na870_1), .IN6(na880_2), .IN7(na850_2),
                      .IN8(na920_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x115y79     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2025_1 ( .OUT(na2025_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na890_2), .IN6(na900_1), .IN7(na910_2),
                      .IN8(na770_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x118y74     80'h00_0018_00_0040_0C0F_5500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2026_1 ( .OUT(na2026_1), .IN1(na2025_1), .IN2(na2024_1), .IN3(na2023_1), .IN4(na2022_1), .IN5(~na2384_1), .IN6(1'b1), .IN7(~na2385_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x128y74     80'h00_0018_00_0040_0C0F_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2027_1 ( .OUT(na2027_1), .IN1(na781_1), .IN2(na861_1), .IN3(na801_2), .IN4(na791_1), .IN5(~na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x130y73     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2028_1 ( .OUT(na2028_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na811_1), .IN6(na821_1), .IN7(na831_1),
                      .IN8(na841_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x125y78     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2029_1 ( .OUT(na2029_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na871_1), .IN6(na881_2), .IN7(na851_2),
                      .IN8(na921_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x127y77     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2030_1 ( .OUT(na2030_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na771_2), .IN6(na911_2), .IN7(na901_1),
                      .IN8(na891_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x126y73     80'h00_0018_00_0040_0C0F_5500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2031_1 ( .OUT(na2031_1), .IN1(na2030_1), .IN2(na2029_1), .IN3(na2028_1), .IN4(na2027_1), .IN5(~na2384_1), .IN6(1'b1), .IN7(~na2385_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x121y32     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2032_1 ( .OUT(na2032_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na932_2), .IN6(na1012_2), .IN7(na952_2),
                      .IN8(na942_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x125y31     80'h00_0018_00_0040_0C0F_5500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2033_1 ( .OUT(na2033_1), .IN1(na992_2), .IN2(na982_2), .IN3(na972_1), .IN4(na962_2), .IN5(~na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x128y32     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2034_1 ( .OUT(na2034_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1002_2), .IN6(na1072_2), .IN7(na1022_2),
                      .IN8(na1032_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x128y31     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2035_1 ( .OUT(na2035_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na922_1), .IN6(na1062_2), .IN7(na1052_2),
                      .IN8(na1042_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x122y29     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2036_1 ( .OUT(na2036_1), .IN1(~na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na2033_1), .IN6(na2032_1), .IN7(na2035_1),
                      .IN8(na2034_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x122y35     80'h00_0018_00_0040_0C0F_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2037_1 ( .OUT(na2037_1), .IN1(na1013_1), .IN2(na933_2), .IN3(na943_1), .IN4(na953_1), .IN5(na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x120y36     80'h00_0018_00_0040_0C0F_5500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2038_1 ( .OUT(na2038_1), .IN1(na993_2), .IN2(na983_2), .IN3(na973_1), .IN4(na963_1), .IN5(~na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x123y39     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2039_1 ( .OUT(na2039_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1003_1), .IN6(na1073_1), .IN7(na1023_1),
                      .IN8(na1033_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x123y38     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2040_1 ( .OUT(na2040_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1043_1), .IN6(na1053_1), .IN7(na1063_2),
                      .IN8(na923_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x124y40     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2041_1 ( .OUT(na2041_1), .IN1(na2384_1), .IN2(1'b1), .IN3(~na2385_1), .IN4(1'b1), .IN5(na2039_1), .IN6(na2040_1), .IN7(na2037_1),
                      .IN8(na2038_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x114y40     80'h00_0018_00_0040_0C0F_5500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2042_1 ( .OUT(na2042_1), .IN1(na954_2), .IN2(na944_1), .IN3(na934_2), .IN4(na1014_1), .IN5(~na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x110y41     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2043_1 ( .OUT(na2043_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na964_2), .IN6(na974_2), .IN7(na984_2),
                      .IN8(na994_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x113y40     80'h00_0018_00_0040_0C0F_5500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2044_1 ( .OUT(na2044_1), .IN1(na1034_2), .IN2(na1024_2), .IN3(na1074_2), .IN4(na1004_2), .IN5(~na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x115y41     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2045_1 ( .OUT(na2045_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1054_2), .IN6(na1044_2), .IN7(na924_2),
                      .IN8(na1064_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x115y42     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2046_1 ( .OUT(na2046_1), .IN1(~na2384_1), .IN2(1'b1), .IN3(~na2385_1), .IN4(1'b1), .IN5(na2045_1), .IN6(na2044_1), .IN7(na2043_1),
                      .IN8(na2042_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x115y45     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2047_1 ( .OUT(na2047_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na955_2), .IN6(na945_1), .IN7(na935_1),
                      .IN8(na1015_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x119y48     80'h00_0018_00_0040_0C0F_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2048_1 ( .OUT(na2048_1), .IN1(na985_1), .IN2(na995_1), .IN3(na965_1), .IN4(na975_1), .IN5(na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x122y49     80'h00_0018_00_0040_0C0F_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2049_1 ( .OUT(na2049_1), .IN1(na1025_1), .IN2(na1035_2), .IN3(na1005_1), .IN4(na1075_1), .IN5(na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x122y48     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2050_1 ( .OUT(na2050_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1055_1), .IN6(na1045_1), .IN7(na925_2),
                      .IN8(na1065_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x117y49     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2051_1 ( .OUT(na2051_1), .IN1(na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na2047_1), .IN6(na2048_1), .IN7(na2049_1),
                      .IN8(na2050_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x112y54     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2052_1 ( .OUT(na2052_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na936_1), .IN6(na1016_2), .IN7(na956_2),
                      .IN8(na946_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x116y53     80'h00_0018_00_0040_0C0F_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2053_1 ( .OUT(na2053_1), .IN1(na986_1), .IN2(na996_2), .IN3(na966_1), .IN4(na976_2), .IN5(na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x113y56     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2054_1 ( .OUT(na2054_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1006_2), .IN6(na1076_2), .IN7(na1026_2),
                      .IN8(na1036_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x115y53     80'h00_0018_00_0040_0C0F_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2055_1 ( .OUT(na2055_1), .IN1(na1056_1), .IN2(na1046_2), .IN3(na926_2), .IN4(na1066_2), .IN5(~na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x115y54     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2056_1 ( .OUT(na2056_1), .IN1(~na2384_1), .IN2(1'b1), .IN3(~na2385_1), .IN4(1'b1), .IN5(na2055_1), .IN6(na2054_1), .IN7(na2053_1),
                      .IN8(na2052_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x117y53     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2057_1 ( .OUT(na2057_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na937_1), .IN6(na1017_1), .IN7(na957_1),
                      .IN8(na947_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x117y54     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2058_1 ( .OUT(na2058_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na997_1), .IN6(na987_1), .IN7(na977_2),
                      .IN8(na967_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x122y55     80'h00_0018_00_0040_0C0F_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2059_1 ( .OUT(na2059_1), .IN1(na1007_2), .IN2(na1077_2), .IN3(na1027_1), .IN4(na1037_1), .IN5(na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x126y54     80'h00_0018_00_0040_0C0F_5500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2060_1 ( .OUT(na2060_1), .IN1(na927_1), .IN2(na1067_1), .IN3(na1057_1), .IN4(na1047_1), .IN5(~na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x120y53     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2061_1 ( .OUT(na2061_1), .IN1(na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na2057_1), .IN6(na2058_1), .IN7(na2059_1),
                      .IN8(na2060_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x118y66     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2062_1 ( .OUT(na2062_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na938_2), .IN6(na1018_2), .IN7(na958_1),
                      .IN8(na948_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x120y65     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2063_1 ( .OUT(na2063_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na998_2), .IN6(na988_2), .IN7(na978_2),
                      .IN8(na968_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x117y66     80'h00_0018_00_0040_0C0F_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2064_1 ( .OUT(na2064_1), .IN1(na1078_2), .IN2(na1008_2), .IN3(na1038_2), .IN4(na1028_1), .IN5(~na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x117y63     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2065_1 ( .OUT(na2065_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1058_2), .IN6(na1048_2), .IN7(na928_1),
                      .IN8(na1068_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x120y62     80'h00_0018_00_0040_0C0F_5500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2066_1 ( .OUT(na2066_1), .IN1(na2065_1), .IN2(na2064_1), .IN3(na2063_1), .IN4(na2062_1), .IN5(~na2384_1), .IN6(1'b1), .IN7(~na2385_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x113y65     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2067_1 ( .OUT(na2067_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na959_1), .IN6(na949_1), .IN7(na939_2),
                      .IN8(na1019_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x115y68     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2068_1 ( .OUT(na2068_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na969_2), .IN6(na979_1), .IN7(na989_1),
                      .IN8(na999_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x114y69     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2069_1 ( .OUT(na2069_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1009_1), .IN6(na1079_1), .IN7(na1029_1),
                      .IN8(na1039_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x116y68     80'h00_0018_00_0040_0C0F_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2070_1 ( .OUT(na2070_1), .IN1(na1069_1), .IN2(na929_1), .IN3(na1049_2), .IN4(na1059_1), .IN5(na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x115y65     80'h00_0018_00_0040_0C0F_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2071_1 ( .OUT(na2071_1), .IN1(na2067_1), .IN2(na2068_1), .IN3(na2069_1), .IN4(na2070_1), .IN5(na2384_1), .IN6(1'b1), .IN7(na2385_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x114y78     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2072_1 ( .OUT(na2072_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na940_2), .IN6(na1020_2), .IN7(na960_2),
                      .IN8(na950_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x116y79     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2073_1 ( .OUT(na2073_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na990_2), .IN6(na1000_1), .IN7(na970_2),
                      .IN8(na980_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x113y74     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2074_1 ( .OUT(na2074_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1010_2), .IN6(na1080_2), .IN7(na1030_2),
                      .IN8(na1040_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x117y79     80'h00_0018_00_0040_0C0F_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2075_1 ( .OUT(na2075_1), .IN1(na1050_2), .IN2(na1060_2), .IN3(na1070_1), .IN4(na930_2), .IN5(na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x118y80     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2076_1 ( .OUT(na2076_1), .IN1(~na2384_1), .IN2(1'b1), .IN3(~na2385_1), .IN4(1'b1), .IN5(na2075_1), .IN6(na2074_1), .IN7(na2073_1),
                      .IN8(na2072_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x136y74     80'h00_0018_00_0040_0C0F_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2077_1 ( .OUT(na2077_1), .IN1(na1021_2), .IN2(na941_1), .IN3(na951_1), .IN4(na961_2), .IN5(na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x136y67     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2078_1 ( .OUT(na2078_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na971_1), .IN6(na981_1), .IN7(na991_1),
                      .IN8(na1001_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x137y70     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2079_1 ( .OUT(na2079_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1081_1), .IN6(na1011_1), .IN7(na1041_1),
                      .IN8(na1031_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x137y67     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2080_1 ( .OUT(na2080_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1061_1), .IN6(na1051_1), .IN7(na931_1),
                      .IN8(na1071_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x135y66     80'h00_0018_00_0040_0C0F_5500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2081_1 ( .OUT(na2081_1), .IN1(na2080_1), .IN2(na2079_1), .IN3(na2078_1), .IN4(na2077_1), .IN5(~na2384_1), .IN6(1'b1), .IN7(~na2385_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x128y36     80'h00_0018_00_0040_0C0F_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2082_1 ( .OUT(na2082_1), .IN1(na1092_2), .IN2(na1172_2), .IN3(na1112_1), .IN4(na1102_2), .IN5(~na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x128y35     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2083_1 ( .OUT(na2083_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1132_2), .IN6(na1122_2), .IN7(na1152_2),
                      .IN8(na1142_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x127y32     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2084_1 ( .OUT(na2084_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1192_2), .IN6(na1182_1), .IN7(na1232_2),
                      .IN8(na1162_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x129y31     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2085_1 ( .OUT(na2085_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1212_2), .IN6(na1202_2), .IN7(na1082_2),
                      .IN8(na1222_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x130y36     80'h00_0018_00_0040_0C0F_5500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2086_1 ( .OUT(na2086_1), .IN1(na2085_1), .IN2(na2084_1), .IN3(na2083_1), .IN4(na2082_1), .IN5(~na2384_1), .IN6(1'b1), .IN7(~na2385_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x125y40     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2087_1 ( .OUT(na2087_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1103_1), .IN6(na1113_1), .IN7(na1173_1),
                      .IN8(na1093_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x129y41     80'h00_0018_00_0040_0C0F_5500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2088_1 ( .OUT(na2088_1), .IN1(na1153_1), .IN2(na1143_1), .IN3(na1133_2), .IN4(na1123_1), .IN5(~na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x130y38     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2089_1 ( .OUT(na2089_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1163_1), .IN6(na1233_1), .IN7(na1183_1),
                      .IN8(na1193_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x130y37     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2090_1 ( .OUT(na2090_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1213_1), .IN6(na1203_2), .IN7(na1083_1),
                      .IN8(na1223_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x127y41     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2091_1 ( .OUT(na2091_1), .IN1(~na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na2088_1), .IN6(na2087_1), .IN7(na2090_1),
                      .IN8(na2089_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x125y39     80'h00_0018_00_0040_0C0F_5500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2092_1 ( .OUT(na2092_1), .IN1(na1114_2), .IN2(na1104_2), .IN3(na1094_2), .IN4(na1174_2), .IN5(~na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x125y34     80'h00_0018_00_0040_0C0F_5500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2093_1 ( .OUT(na2093_1), .IN1(na1154_1), .IN2(na1144_2), .IN3(na1134_2), .IN4(na1124_2), .IN5(~na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x124y35     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2094_1 ( .OUT(na2094_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1184_2), .IN6(na1194_2), .IN7(na1164_2),
                      .IN8(na1234_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x124y38     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2095_1 ( .OUT(na2095_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1214_2), .IN6(na1204_2), .IN7(na1084_1),
                      .IN8(na1224_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x125y41     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2096_1 ( .OUT(na2096_1), .IN1(na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na2092_1), .IN6(na2093_1), .IN7(na2094_1),
                      .IN8(na2095_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x134y44     80'h00_0018_00_0040_0C0F_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2097_1 ( .OUT(na2097_1), .IN1(na1105_2), .IN2(na1115_1), .IN3(na1175_2), .IN4(na1095_1), .IN5(na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x136y47     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2098_1 ( .OUT(na2098_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1125_1), .IN6(na1135_1), .IN7(na1145_1),
                      .IN8(na1155_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x129y48     80'h00_0018_00_0040_0C0F_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2099_1 ( .OUT(na2099_1), .IN1(na1235_1), .IN2(na1165_1), .IN3(na1195_1), .IN4(na1185_1), .IN5(~na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x131y45     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2100_1 ( .OUT(na2100_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1205_1), .IN6(na1215_1), .IN7(na1225_1),
                      .IN8(na1085_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x137y51     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2101_1 ( .OUT(na2101_1), .IN1(~na2384_1), .IN2(1'b1), .IN3(~na2385_1), .IN4(1'b1), .IN5(na2100_1), .IN6(na2099_1), .IN7(na2098_1),
                      .IN8(na2097_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x134y56     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2102_1 ( .OUT(na2102_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1176_2), .IN6(na1096_2), .IN7(na1106_2),
                      .IN8(na1116_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x134y55     80'h00_0018_00_0040_0C0F_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2103_1 ( .OUT(na2103_1), .IN1(na1146_2), .IN2(na1156_2), .IN3(na1126_1), .IN4(na1136_2), .IN5(na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x133y56     80'h00_0018_00_0040_0C0F_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2104_1 ( .OUT(na2104_1), .IN1(na1186_2), .IN2(na1196_1), .IN3(na1166_2), .IN4(na1236_2), .IN5(na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x135y55     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2105_1 ( .OUT(na2105_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1086_2), .IN6(na1226_2), .IN7(na1216_2),
                      .IN8(na1206_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x133y55     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2106_1 ( .OUT(na2106_1), .IN1(~na2384_1), .IN2(1'b1), .IN3(~na2385_1), .IN4(1'b1), .IN5(na2105_1), .IN6(na2104_1), .IN7(na2103_1),
                      .IN8(na2102_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x123y63     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2107_1 ( .OUT(na2107_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1107_1), .IN6(na1117_1), .IN7(na1177_1),
                      .IN8(na1097_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x123y64     80'h00_0018_00_0040_0C0F_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2108_1 ( .OUT(na2108_1), .IN1(na1127_1), .IN2(na1137_1), .IN3(na1147_2), .IN4(na1157_1), .IN5(na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x124y61     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2109_1 ( .OUT(na2109_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1187_1), .IN6(na1197_1), .IN7(na1167_1),
                      .IN8(na1237_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x122y60     80'h00_0018_00_0040_0C0F_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2110_1 ( .OUT(na2110_1), .IN1(na1227_1), .IN2(na1087_1), .IN3(na1207_1), .IN4(na1217_2), .IN5(na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x123y59     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2111_1 ( .OUT(na2111_1), .IN1(na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na2107_1), .IN6(na2108_1), .IN7(na2109_1),
                      .IN8(na2110_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x117y69     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2112_1 ( .OUT(na2112_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1098_1), .IN6(na1178_2), .IN7(na1118_2),
                      .IN8(na1108_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x119y70     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2113_1 ( .OUT(na2113_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1158_2), .IN6(na1148_2), .IN7(na1138_2),
                      .IN8(na1128_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x122y67     80'h00_0018_00_0040_0C0F_5500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2114_1 ( .OUT(na2114_1), .IN1(na1198_2), .IN2(na1188_2), .IN3(na1238_1), .IN4(na1168_1), .IN5(~na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x118y68     80'h00_0018_00_0040_0C0F_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2115_1 ( .OUT(na2115_1), .IN1(na1228_2), .IN2(na1088_2), .IN3(na1208_2), .IN4(na1218_2), .IN5(na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x118y63     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2116_1 ( .OUT(na2116_1), .IN1(na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na2112_1), .IN6(na2113_1), .IN7(na2114_1),
                      .IN8(na2115_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x118y69     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2117_1 ( .OUT(na2117_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1179_1), .IN6(na1099_1), .IN7(na1109_1),
                      .IN8(na1119_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x120y74     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2118_1 ( .OUT(na2118_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1129_1), .IN6(na1139_1), .IN7(na1149_1),
                      .IN8(na1159_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x119y69     80'h00_0018_00_0040_0C0F_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2119_1 ( .OUT(na2119_1), .IN1(na1189_2), .IN2(na1199_1), .IN3(na1169_1), .IN4(na1239_1), .IN5(na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x119y76     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2120_1 ( .OUT(na2120_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1229_1), .IN6(na1089_1), .IN7(na1209_1),
                      .IN8(na1219_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x118y67     80'h00_0018_00_0040_0C0F_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2121_1 ( .OUT(na2121_1), .IN1(na2119_1), .IN2(na2120_1), .IN3(na2117_1), .IN4(na2118_1), .IN5(na2384_1), .IN6(1'b1), .IN7(~na2385_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x127y72     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2122_1 ( .OUT(na2122_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1180_2), .IN6(na1100_2), .IN7(na1110_2),
                      .IN8(na1120_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x129y71     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2123_1 ( .OUT(na2123_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1150_2), .IN6(na1160_2), .IN7(na1130_2),
                      .IN8(na1140_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x130y72     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2124_1 ( .OUT(na2124_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1170_2), .IN6(na1240_2), .IN7(na1190_2),
                      .IN8(na1200_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x130y75     80'h00_0018_00_0040_0C0F_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2125_1 ( .OUT(na2125_1), .IN1(na1210_1), .IN2(na1220_2), .IN3(na1230_2), .IN4(na1090_2), .IN5(na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x128y70     80'h00_0018_00_0040_0C0F_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2126_1 ( .OUT(na2126_1), .IN1(na2123_1), .IN2(na2122_1), .IN3(na2125_1), .IN4(na2124_1), .IN5(~na2384_1), .IN6(1'b1), .IN7(na2385_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x131y77     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2127_1 ( .OUT(na2127_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1101_1), .IN6(na1181_1), .IN7(na1121_1),
                      .IN8(na1111_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x129y82     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2128_1 ( .OUT(na2128_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1141_1), .IN6(na1131_1), .IN7(na1161_2),
                      .IN8(na1151_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x132y75     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2129_1 ( .OUT(na2129_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1171_1), .IN6(na1241_1), .IN7(na1191_1),
                      .IN8(na1201_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x128y84     80'h00_0018_00_0040_0C0F_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2130_1 ( .OUT(na2130_1), .IN1(na1231_2), .IN2(na1091_2), .IN3(na1211_1), .IN4(na1221_1), .IN5(na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x130y77     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2131_1 ( .OUT(na2131_1), .IN1(na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na2127_1), .IN6(na2128_1), .IN7(na2129_1),
                      .IN8(na2130_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x153y37     80'h00_0018_00_0040_0C0F_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2132_1 ( .OUT(na2132_1), .IN1(na1252_1), .IN2(na1332_2), .IN3(na1272_2), .IN4(na1262_2), .IN5(~na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x151y36     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2133_1 ( .OUT(na2133_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1292_2), .IN6(na1282_2), .IN7(na1312_2),
                      .IN8(na1302_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x152y39     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2134_1 ( .OUT(na2134_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1342_2), .IN6(na1352_2), .IN7(na1322_1),
                      .IN8(na1392_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x152y36     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2135_1 ( .OUT(na2135_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1382_2), .IN6(na1242_2), .IN7(na1362_2),
                      .IN8(na1372_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x148y42     80'h00_0018_00_0040_0C0F_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2136_1 ( .OUT(na2136_1), .IN1(na2132_1), .IN2(na2133_1), .IN3(na2134_1), .IN4(na2135_1), .IN5(na2384_1), .IN6(1'b1), .IN7(na2385_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x130y41     80'h00_0018_00_0040_0C0F_5500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2137_1 ( .OUT(na2137_1), .IN1(na1273_2), .IN2(na1263_1), .IN3(na1253_1), .IN4(na1333_1), .IN5(~na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x130y40     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2138_1 ( .OUT(na2138_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1313_1), .IN6(na1303_1), .IN7(na1293_1),
                      .IN8(na1283_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x129y45     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2139_1 ( .OUT(na2139_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1353_1), .IN6(na1343_2), .IN7(na1393_1),
                      .IN8(na1323_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x133y38     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2140_1 ( .OUT(na2140_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1243_1), .IN6(na1383_1), .IN7(na1373_1),
                      .IN8(na1363_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x134y42     80'h00_0018_00_0040_0C0F_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2141_1 ( .OUT(na2141_1), .IN1(na2139_1), .IN2(na2140_1), .IN3(na2137_1), .IN4(na2138_1), .IN5(na2384_1), .IN6(1'b1), .IN7(~na2385_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x152y44     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2142_1 ( .OUT(na2142_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1264_2), .IN6(na1274_2), .IN7(na1334_2),
                      .IN8(na1254_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x150y43     80'h00_0018_00_0040_0C0F_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2143_1 ( .OUT(na2143_1), .IN1(na1304_2), .IN2(na1314_2), .IN3(na1284_2), .IN4(na1294_1), .IN5(na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x149y44     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2144_1 ( .OUT(na2144_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1324_2), .IN6(na1394_2), .IN7(na1344_2),
                      .IN8(na1354_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x149y45     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2145_1 ( .OUT(na2145_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1384_2), .IN6(na1244_2), .IN7(na1364_1),
                      .IN8(na1374_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x150y46     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2146_1 ( .OUT(na2146_1), .IN1(~na2384_1), .IN2(1'b1), .IN3(~na2385_1), .IN4(1'b1), .IN5(na2145_1), .IN6(na2144_1), .IN7(na2143_1),
                      .IN8(na2142_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x133y53     80'h00_0018_00_0040_0C0F_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2147_1 ( .OUT(na2147_1), .IN1(na1265_1), .IN2(na1275_1), .IN3(na1335_1), .IN4(na1255_1), .IN5(na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x137y54     80'h00_0018_00_0040_0C0F_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2148_1 ( .OUT(na2148_1), .IN1(na1295_1), .IN2(na1285_1), .IN3(na1315_2), .IN4(na1305_1), .IN5(~na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x138y51     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2149_1 ( .OUT(na2149_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1325_1), .IN6(na1395_1), .IN7(na1345_1),
                      .IN8(na1355_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x140y52     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2150_1 ( .OUT(na2150_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1375_1), .IN6(na1365_1), .IN7(na1245_2),
                      .IN8(na1385_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x138y52     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2151_1 ( .OUT(na2151_1), .IN1(na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na2147_1), .IN6(na2148_1), .IN7(na2149_1),
                      .IN8(na2150_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x151y50     80'h00_0018_00_0040_0C0F_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2152_1 ( .OUT(na2152_1), .IN1(na1256_2), .IN2(na1336_1), .IN3(na1276_2), .IN4(na1266_1), .IN5(~na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x151y49     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2153_1 ( .OUT(na2153_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1306_2), .IN6(na1316_2), .IN7(na1286_2),
                      .IN8(na1296_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x154y48     80'h00_0018_00_0040_0C0F_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2154_1 ( .OUT(na2154_1), .IN1(na1346_2), .IN2(na1356_2), .IN3(na1326_2), .IN4(na1396_2), .IN5(na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x154y45     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2155_1 ( .OUT(na2155_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1366_2), .IN6(na1376_2), .IN7(na1386_2),
                      .IN8(na1246_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x148y50     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2156_1 ( .OUT(na2156_1), .IN1(~na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na2153_1), .IN6(na2152_1), .IN7(na2155_1),
                      .IN8(na2154_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x151y56     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2157_1 ( .OUT(na2157_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1277_1), .IN6(na1267_1), .IN7(na1257_1),
                      .IN8(na1337_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x151y55     80'h00_0018_00_0040_0C0F_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2158_1 ( .OUT(na2158_1), .IN1(na1287_2), .IN2(na1297_1), .IN3(na1307_1), .IN4(na1317_1), .IN5(na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x154y58     80'h00_0018_00_0040_0C0F_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2159_1 ( .OUT(na2159_1), .IN1(na1347_1), .IN2(na1357_2), .IN3(na1327_1), .IN4(na1397_1), .IN5(na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x152y55     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2160_1 ( .OUT(na2160_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1367_1), .IN6(na1377_1), .IN7(na1387_1),
                      .IN8(na1247_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x148y58     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2161_1 ( .OUT(na2161_1), .IN1(~na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na2158_1), .IN6(na2157_1), .IN7(na2160_1),
                      .IN8(na2159_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x144y68     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2162_1 ( .OUT(na2162_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1268_2), .IN6(na1278_2), .IN7(na1338_2),
                      .IN8(na1258_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x150y65     80'h00_0018_00_0040_0C0F_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2163_1 ( .OUT(na2163_1), .IN1(na1298_2), .IN2(na1288_2), .IN3(na1318_2), .IN4(na1308_1), .IN5(~na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x147y68     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2164_1 ( .OUT(na2164_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1398_2), .IN6(na1328_2), .IN7(na1358_2),
                      .IN8(na1348_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x145y69     80'h00_0018_00_0040_0C0F_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2165_1 ( .OUT(na2165_1), .IN1(na1388_2), .IN2(na1248_2), .IN3(na1368_2), .IN4(na1378_1), .IN5(na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x144y66     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2166_1 ( .OUT(na2166_1), .IN1(~na2384_1), .IN2(1'b1), .IN3(~na2385_1), .IN4(1'b1), .IN5(na2165_1), .IN6(na2164_1), .IN7(na2163_1),
                      .IN8(na2162_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x151y73     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2167_1 ( .OUT(na2167_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1339_1), .IN6(na1259_2), .IN7(na1269_1),
                      .IN8(na1279_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x145y72     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2168_1 ( .OUT(na2168_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1309_1), .IN6(na1319_1), .IN7(na1289_1),
                      .IN8(na1299_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x148y69     80'h00_0018_00_0040_0C0F_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2169_1 ( .OUT(na2169_1), .IN1(na1329_2), .IN2(na1399_2), .IN3(na1349_1), .IN4(na1359_1), .IN5(na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x152y72     80'h00_0018_00_0040_0C0F_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2170_1 ( .OUT(na2170_1), .IN1(na1379_1), .IN2(na1369_1), .IN3(na1249_1), .IN4(na1389_1), .IN5(~na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x152y70     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2171_1 ( .OUT(na2171_1), .IN1(na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na2167_1), .IN6(na2168_1), .IN7(na2169_1),
                      .IN8(na2170_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x153y77     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2172_1 ( .OUT(na2172_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1340_2), .IN6(na1260_2), .IN7(na1270_2),
                      .IN8(na1280_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x153y80     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2173_1 ( .OUT(na2173_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1320_2), .IN6(na1310_2), .IN7(na1300_2),
                      .IN8(na1290_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x152y75     80'h00_0018_00_0040_0C0F_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2174_1 ( .OUT(na2174_1), .IN1(na1330_2), .IN2(na1400_2), .IN3(na1350_1), .IN4(na1360_2), .IN5(na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x152y80     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2175_1 ( .OUT(na2175_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1380_2), .IN6(na1370_2), .IN7(na1250_2),
                      .IN8(na1390_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x152y76     80'h00_0018_00_0040_0C0F_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2176_1 ( .OUT(na2176_1), .IN1(na2172_1), .IN2(na2173_1), .IN3(na2174_1), .IN4(na2175_1), .IN5(na2384_1), .IN6(1'b1), .IN7(na2385_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x145y80     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2177_1 ( .OUT(na2177_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1281_1), .IN6(na1271_1), .IN7(na1261_1),
                      .IN8(na1341_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x141y75     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2178_1 ( .OUT(na2178_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1291_1), .IN6(na1301_2), .IN7(na1311_1),
                      .IN8(na1321_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x142y76     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2179_1 ( .OUT(na2179_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1351_1), .IN6(na1361_1), .IN7(na1331_1),
                      .IN8(na1401_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x142y81     80'h00_0018_00_0040_0C0F_5500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2180_1 ( .OUT(na2180_1), .IN1(na1251_1), .IN2(na1391_1), .IN3(na1381_1), .IN4(na1371_2), .IN5(~na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x144y76     80'h00_0018_00_0040_0C0F_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2181_1 ( .OUT(na2181_1), .IN1(na2178_1), .IN2(na2177_1), .IN3(na2180_1), .IN4(na2179_1), .IN5(~na2384_1), .IN6(1'b1), .IN7(na2385_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x112y33     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2182_1 ( .OUT(na2182_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1492_2), .IN6(na1412_2), .IN7(na1422_2),
                      .IN8(na1432_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x116y34     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2183_1 ( .OUT(na2183_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1452_2), .IN6(na1442_2), .IN7(na1472_2),
                      .IN8(na1462_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x115y33     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2184_1 ( .OUT(na2184_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1512_2), .IN6(na1502_2), .IN7(na1552_2),
                      .IN8(na1482_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x117y36     80'h00_0018_00_0040_0C0F_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2185_1 ( .OUT(na2185_1), .IN1(na1522_2), .IN2(na1532_1), .IN3(na1542_2), .IN4(na1402_2), .IN5(na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x115y34     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2186_1 ( .OUT(na2186_1), .IN1(na2384_1), .IN2(1'b1), .IN3(~na2385_1), .IN4(1'b1), .IN5(na2184_1), .IN6(na2185_1), .IN7(na2182_1),
                      .IN8(na2183_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x111y33     80'h00_0018_00_0040_0C0F_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2187_1 ( .OUT(na2187_1), .IN1(na1413_2), .IN2(na1493_1), .IN3(na1433_1), .IN4(na1423_1), .IN5(~na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x115y38     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2188_1 ( .OUT(na2188_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1453_1), .IN6(na1443_1), .IN7(na1473_1),
                      .IN8(na1463_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x116y35     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2189_1 ( .OUT(na2189_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1513_1), .IN6(na1503_1), .IN7(na1553_2),
                      .IN8(na1483_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x114y36     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2190_1 ( .OUT(na2190_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1523_1), .IN6(na1533_1), .IN7(na1543_1),
                      .IN8(na1403_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x112y39     80'h00_0018_00_0040_0C0F_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2191_1 ( .OUT(na2191_1), .IN1(na2187_1), .IN2(na2188_1), .IN3(na2189_1), .IN4(na2190_1), .IN5(na2384_1), .IN6(1'b1), .IN7(na2385_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x110y39     80'h00_0018_00_0040_0C0F_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2192_1 ( .OUT(na2192_1), .IN1(na1424_2), .IN2(na1434_1), .IN3(na1494_2), .IN4(na1414_2), .IN5(na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x110y40     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2193_1 ( .OUT(na2193_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1454_2), .IN6(na1444_2), .IN7(na1474_2),
                      .IN8(na1464_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x113y43     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2194_1 ( .OUT(na2194_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1484_2), .IN6(na1554_2), .IN7(na1504_1),
                      .IN8(na1514_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x107y42     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2195_1 ( .OUT(na2195_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1534_2), .IN6(na1524_2), .IN7(na1404_2),
                      .IN8(na1544_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x111y42     80'h00_0018_00_0040_0C0F_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2196_1 ( .OUT(na2196_1), .IN1(na2194_1), .IN2(na2195_1), .IN3(na2192_1), .IN4(na2193_1), .IN5(na2384_1), .IN6(1'b1), .IN7(~na2385_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x110y46     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2197_1 ( .OUT(na2197_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1425_1), .IN6(na1435_1), .IN7(na1495_1),
                      .IN8(na1415_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x112y47     80'h00_0018_00_0040_0C0F_5500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2198_1 ( .OUT(na2198_1), .IN1(na1475_1), .IN2(na1465_1), .IN3(na1455_2), .IN4(na1445_1), .IN5(~na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x113y44     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2199_1 ( .OUT(na2199_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1485_1), .IN6(na1555_1), .IN7(na1505_1),
                      .IN8(na1515_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x109y47     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2200_1 ( .OUT(na2200_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1525_2), .IN6(na1535_1), .IN7(na1545_1),
                      .IN8(na1405_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x113y45     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2201_1 ( .OUT(na2201_1), .IN1(~na2384_1), .IN2(1'b1), .IN3(~na2385_1), .IN4(1'b1), .IN5(na2200_1), .IN6(na2199_1), .IN7(na2198_1),
                      .IN8(na2197_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x106y58     80'h00_0018_00_0040_0C0F_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2202_1 ( .OUT(na2202_1), .IN1(na1416_2), .IN2(na1496_2), .IN3(na1436_2), .IN4(na1426_2), .IN5(~na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x110y59     80'h00_0018_00_0040_0C0F_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2203_1 ( .OUT(na2203_1), .IN1(na1466_2), .IN2(na1476_1), .IN3(na1446_2), .IN4(na1456_2), .IN5(na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x107y58     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2204_1 ( .OUT(na2204_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1516_2), .IN6(na1506_2), .IN7(na1556_2),
                      .IN8(na1486_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x111y59     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2205_1 ( .OUT(na2205_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1406_1), .IN6(na1546_1), .IN7(na1536_2),
                      .IN8(na1526_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x108y58     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2206_1 ( .OUT(na2206_1), .IN1(~na2384_1), .IN2(1'b1), .IN3(~na2385_1), .IN4(1'b1), .IN5(na2205_1), .IN6(na2204_1), .IN7(na2203_1),
                      .IN8(na2202_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x115y61     80'h00_0018_00_0040_0C0F_5500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2207_1 ( .OUT(na2207_1), .IN1(na1437_1), .IN2(na1427_2), .IN3(na1417_1), .IN4(na1497_2), .IN5(~na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x119y62     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2208_1 ( .OUT(na2208_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1447_1), .IN6(na1457_1), .IN7(na1467_1),
                      .IN8(na1477_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x120y61     80'h00_0018_00_0040_0C0F_5500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2209_1 ( .OUT(na2209_1), .IN1(na1517_1), .IN2(na1507_1), .IN3(na1557_1), .IN4(na1487_1), .IN5(~na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x118y62     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2210_1 ( .OUT(na2210_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1547_1), .IN6(na1407_1), .IN7(na1527_1),
                      .IN8(na1537_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x120y60     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2211_1 ( .OUT(na2211_1), .IN1(na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na2207_1), .IN6(na2208_1), .IN7(na2209_1),
                      .IN8(na2210_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x105y64     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2212_1 ( .OUT(na2212_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1498_2), .IN6(na1418_2), .IN7(na1428_2),
                      .IN8(na1438_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x107y65     80'h00_0018_00_0040_0C0F_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2213_1 ( .OUT(na2213_1), .IN1(na1468_2), .IN2(na1478_2), .IN3(na1448_1), .IN4(na1458_2), .IN5(na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x110y66     80'h00_0018_00_0040_0C0F_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2214_1 ( .OUT(na2214_1), .IN1(na1508_2), .IN2(na1518_1), .IN3(na1488_2), .IN4(na1558_2), .IN5(na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x106y67     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2215_1 ( .OUT(na2215_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1538_2), .IN6(na1528_2), .IN7(na1408_2),
                      .IN8(na1548_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x112y64     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2216_1 ( .OUT(na2216_1), .IN1(~na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na2213_1), .IN6(na2212_1), .IN7(na2215_1),
                      .IN8(na2214_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x111y69     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2217_1 ( .OUT(na2217_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1429_1), .IN6(na1439_1), .IN7(na1499_1),
                      .IN8(na1419_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x111y74     80'h00_0018_00_0040_0C0F_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2218_1 ( .OUT(na2218_1), .IN1(na1449_1), .IN2(na1459_1), .IN3(na1469_2), .IN4(na1479_1), .IN5(na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x112y73     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2219_1 ( .OUT(na2219_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1559_1), .IN6(na1489_1), .IN7(na1519_1),
                      .IN8(na1509_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x110y76     80'h00_0018_00_0040_0C0F_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2220_1 ( .OUT(na2220_1), .IN1(na1529_1), .IN2(na1539_2), .IN3(na1549_1), .IN4(na1409_1), .IN5(na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x115y69     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2221_1 ( .OUT(na2221_1), .IN1(na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na2217_1), .IN6(na2218_1), .IN7(na2219_1),
                      .IN8(na2220_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x109y82     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2222_1 ( .OUT(na2222_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1500_2), .IN6(na1420_1), .IN7(na1430_2),
                      .IN8(na1440_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x111y81     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2223_1 ( .OUT(na2223_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1470_2), .IN6(na1480_2), .IN7(na1450_2),
                      .IN8(na1460_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x116y84     80'h00_0018_00_0040_0C0F_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2224_1 ( .OUT(na2224_1), .IN1(na1510_2), .IN2(na1520_2), .IN3(na1490_1), .IN4(na1560_1), .IN5(na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x112y81     80'h00_0018_00_0040_0C0F_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2225_1 ( .OUT(na2225_1), .IN1(na1530_2), .IN2(na1540_2), .IN3(na1550_2), .IN4(na1410_2), .IN5(na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x115y81     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2226_1 ( .OUT(na2226_1), .IN1(~na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na2223_1), .IN6(na2222_1), .IN7(na2225_1),
                      .IN8(na2224_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x124y81     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2227_1 ( .OUT(na2227_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1441_2), .IN6(na1431_1), .IN7(na1421_1),
                      .IN8(na1501_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x124y76     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2228_1 ( .OUT(na2228_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1461_1), .IN6(na1451_1), .IN7(na1481_1),
                      .IN8(na1471_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x123y75     80'h00_0018_00_0040_0C0F_5500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2229_1 ( .OUT(na2229_1), .IN1(na1521_1), .IN2(na1511_2), .IN3(na1561_1), .IN4(na1491_1), .IN5(~na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x123y78     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2230_1 ( .OUT(na2230_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1411_1), .IN6(na1551_1), .IN7(na1541_1),
                      .IN8(na1531_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x123y72     80'h00_0018_00_0040_0C0F_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2231_1 ( .OUT(na2231_1), .IN1(na2229_1), .IN2(na2230_1), .IN3(na2227_1), .IN4(na2228_1), .IN5(na2384_1), .IN6(1'b1), .IN7(~na2385_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x132y31     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2232_1 ( .OUT(na2232_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1572_2), .IN6(na1652_2), .IN7(na1592_2),
                      .IN8(na1582_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x134y32     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2233_1 ( .OUT(na2233_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1622_2), .IN6(na1632_2), .IN7(na1602_1),
                      .IN8(na1612_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x131y31     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2234_1 ( .OUT(na2234_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1642_2), .IN6(na1712_2), .IN7(na1662_2),
                      .IN8(na1672_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x135y32     80'h00_0018_00_0040_0C0F_5500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2235_1 ( .OUT(na2235_1), .IN1(na1562_2), .IN2(na1702_2), .IN3(na1692_2), .IN4(na1682_2), .IN5(~na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x131y34     80'h00_0018_00_0040_0C0F_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2236_1 ( .OUT(na2236_1), .IN1(na2234_1), .IN2(na2235_1), .IN3(na2232_1), .IN4(na2233_1), .IN5(na2384_1), .IN6(1'b1), .IN7(~na2385_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x133y35     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2237_1 ( .OUT(na2237_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1593_1), .IN6(na1583_1), .IN7(na1573_1),
                      .IN8(na1653_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x135y36     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2238_1 ( .OUT(na2238_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1603_1), .IN6(na1613_1), .IN7(na1623_2),
                      .IN8(na1633_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x136y35     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2239_1 ( .OUT(na2239_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1673_1), .IN6(na1663_1), .IN7(na1713_1),
                      .IN8(na1643_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x136y34     80'h00_0018_00_0040_0C0F_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2240_1 ( .OUT(na2240_1), .IN1(na1683_1), .IN2(na1693_2), .IN3(na1703_1), .IN4(na1563_1), .IN5(na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x137y37     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2241_1 ( .OUT(na2241_1), .IN1(na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na2237_1), .IN6(na2238_1), .IN7(na2239_1),
                      .IN8(na2240_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x127y44     80'h00_0018_00_0040_0C0F_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2242_1 ( .OUT(na2242_1), .IN1(na1574_1), .IN2(na1654_2), .IN3(na1594_2), .IN4(na1584_2), .IN5(~na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x127y47     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2243_1 ( .OUT(na2243_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1634_2), .IN6(na1624_2), .IN7(na1614_2),
                      .IN8(na1604_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x128y44     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2244_1 ( .OUT(na2244_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1674_2), .IN6(na1664_2), .IN7(na1714_1),
                      .IN8(na1644_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x128y41     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2245_1 ( .OUT(na2245_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1684_2), .IN6(na1694_2), .IN7(na1704_2),
                      .IN8(na1564_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x126y44     80'h00_0018_00_0040_0C0F_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2246_1 ( .OUT(na2246_1), .IN1(na2243_1), .IN2(na2242_1), .IN3(na2245_1), .IN4(na2244_1), .IN5(~na2384_1), .IN6(1'b1), .IN7(na2385_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x140y46     80'h00_0018_00_0040_0C0F_5500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2247_1 ( .OUT(na2247_1), .IN1(na1595_2), .IN2(na1585_1), .IN3(na1575_1), .IN4(na1655_1), .IN5(~na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x140y45     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2248_1 ( .OUT(na2248_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1625_1), .IN6(na1635_1), .IN7(na1605_1),
                      .IN8(na1615_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x139y46     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2249_1 ( .OUT(na2249_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1675_1), .IN6(na1665_2), .IN7(na1715_1),
                      .IN8(na1645_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x141y45     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2250_1 ( .OUT(na2250_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1565_1), .IN6(na1705_1), .IN7(na1695_1),
                      .IN8(na1685_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x141y43     80'h00_0018_00_0040_0C0F_5500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2251_1 ( .OUT(na2251_1), .IN1(na2250_1), .IN2(na2249_1), .IN3(na2248_1), .IN4(na2247_1), .IN5(~na2384_1), .IN6(1'b1), .IN7(~na2385_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x131y62     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2252_1 ( .OUT(na2252_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1576_2), .IN6(na1656_2), .IN7(na1596_2),
                      .IN8(na1586_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x129y63     80'h00_0018_00_0040_0C0F_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2253_1 ( .OUT(na2253_1), .IN1(na1616_1), .IN2(na1606_2), .IN3(na1636_2), .IN4(na1626_2), .IN5(~na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x134y64     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2254_1 ( .OUT(na2254_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1646_2), .IN6(na1716_2), .IN7(na1666_2),
                      .IN8(na1676_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x132y63     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2255_1 ( .OUT(na2255_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1566_2), .IN6(na1706_2), .IN7(na1696_2),
                      .IN8(na1686_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x131y61     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2256_1 ( .OUT(na2256_1), .IN1(~na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na2253_1), .IN6(na2252_1), .IN7(na2255_1),
                      .IN8(na2254_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x138y59     80'h00_0018_00_0040_0C0F_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2257_1 ( .OUT(na2257_1), .IN1(na1657_1), .IN2(na1577_1), .IN3(na1587_1), .IN4(na1597_1), .IN5(na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x138y62     80'h00_0018_00_0040_0C0F_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2258_1 ( .OUT(na2258_1), .IN1(na1607_1), .IN2(na1617_1), .IN3(na1627_1), .IN4(na1637_2), .IN5(na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x137y65     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2259_1 ( .OUT(na2259_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1677_1), .IN6(na1667_1), .IN7(na1717_1),
                      .IN8(na1647_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x139y64     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2260_1 ( .OUT(na2260_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1707_2), .IN6(na1567_2), .IN7(na1687_1),
                      .IN8(na1697_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x140y59     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2261_1 ( .OUT(na2261_1), .IN1(na2384_1), .IN2(1'b1), .IN3(~na2385_1), .IN4(1'b1), .IN5(na2259_1), .IN6(na2260_1), .IN7(na2257_1),
                      .IN8(na2258_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x126y70     80'h00_0018_00_0040_0C0F_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2262_1 ( .OUT(na2262_1), .IN1(na1588_1), .IN2(na1598_2), .IN3(na1658_1), .IN4(na1578_2), .IN5(na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x130y69     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2263_1 ( .OUT(na2263_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1608_2), .IN6(na1618_2), .IN7(na1628_2),
                      .IN8(na1638_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x129y72     80'h00_0018_00_0040_0C0F_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2264_1 ( .OUT(na2264_1), .IN1(na1718_2), .IN2(na1648_2), .IN3(na1678_2), .IN4(na1668_2), .IN5(~na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x131y69     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2265_1 ( .OUT(na2265_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1698_2), .IN6(na1688_2), .IN7(na1568_2),
                      .IN8(na1708_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x124y68     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2266_1 ( .OUT(na2266_1), .IN1(~na2384_1), .IN2(1'b1), .IN3(~na2385_1), .IN4(1'b1), .IN5(na2265_1), .IN6(na2264_1), .IN7(na2263_1),
                      .IN8(na2262_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x133y67     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2267_1 ( .OUT(na2267_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1599_1), .IN6(na1589_1), .IN7(na1579_1),
                      .IN8(na1659_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x133y68     80'h00_0018_00_0040_0C0F_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2268_1 ( .OUT(na2268_1), .IN1(na1629_1), .IN2(na1639_1), .IN3(na1609_2), .IN4(na1619_1), .IN5(na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x130y71     80'h00_0018_00_0040_0C0F_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2269_1 ( .OUT(na2269_1), .IN1(na1669_1), .IN2(na1679_2), .IN3(na1649_1), .IN4(na1719_1), .IN5(na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x132y72     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2270_1 ( .OUT(na2270_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1569_1), .IN6(na1709_1), .IN7(na1699_1),
                      .IN8(na1689_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x135y67     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2271_1 ( .OUT(na2271_1), .IN1(na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na2267_1), .IN6(na2268_1), .IN7(na2269_1),
                      .IN8(na2270_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x131y73     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2272_1 ( .OUT(na2272_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1580_2), .IN6(na1660_2), .IN7(na1600_2),
                      .IN8(na1590_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x133y74     80'h00_0018_00_0040_0C0F_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2273_1 ( .OUT(na2273_1), .IN1(na1610_2), .IN2(na1620_2), .IN3(na1630_1), .IN4(na1640_2), .IN5(na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x138y75     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2274_1 ( .OUT(na2274_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1670_2), .IN6(na1680_2), .IN7(na1650_2),
                      .IN8(na1720_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x134y76     80'h00_0018_00_0040_0C0F_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2275_1 ( .OUT(na2275_1), .IN1(na1700_1), .IN2(na1690_2), .IN3(na1570_2), .IN4(na1710_2), .IN5(~na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x133y72     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2276_1 ( .OUT(na2276_1), .IN1(na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na2272_1), .IN6(na2273_1), .IN7(na2274_1),
                      .IN8(na2275_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x145y81     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2277_1 ( .OUT(na2277_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1661_1), .IN6(na1581_2), .IN7(na1591_1),
                      .IN8(na1601_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x145y82     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2278_1 ( .OUT(na2278_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1611_1), .IN6(na1621_1), .IN7(na1631_1),
                      .IN8(na1641_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x152y79     80'h00_0018_00_0040_0C0F_5500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2279_1 ( .OUT(na2279_1), .IN1(na1681_1), .IN2(na1671_1), .IN3(na1721_2), .IN4(na1651_2), .IN5(~na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x148y82     80'h00_0018_00_0040_0C0F_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2280_1 ( .OUT(na2280_1), .IN1(na1691_1), .IN2(na1701_1), .IN3(na1711_1), .IN4(na1571_1), .IN5(na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x147y79     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2281_1 ( .OUT(na2281_1), .IN1(na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na2277_1), .IN6(na2278_1), .IN7(na2279_1),
                      .IN8(na2280_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x155y36     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2282_1 ( .OUT(na2282_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1812_1), .IN6(na1732_2), .IN7(na1742_1),
                      .IN8(na1752_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x153y33     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2283_1 ( .OUT(na2283_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1762_2), .IN6(na1772_2), .IN7(na1782_2),
                      .IN8(na1792_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x152y32     80'h00_0018_00_0040_0C0F_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2284_1 ( .OUT(na2284_1), .IN1(na1822_2), .IN2(na1832_2), .IN3(na1802_2), .IN4(na1872_2), .IN5(na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x154y33     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2285_1 ( .OUT(na2285_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1842_2), .IN6(na1852_2), .IN7(na1862_2),
                      .IN8(na1722_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x154y36     80'h00_0018_00_0040_0C0F_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2286_1 ( .OUT(na2286_1), .IN1(na2283_1), .IN2(na2282_1), .IN3(na2285_1), .IN4(na2284_1), .IN5(~na2384_1), .IN6(1'b1), .IN7(na2385_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x135y41     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2287_1 ( .OUT(na2287_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1813_1), .IN6(na1733_1), .IN7(na1743_1),
                      .IN8(na1753_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x139y40     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2288_1 ( .OUT(na2288_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1763_2), .IN6(na1773_1), .IN7(na1783_1),
                      .IN8(na1793_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x142y39     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2289_1 ( .OUT(na2289_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1823_1), .IN6(na1833_2), .IN7(na1803_1),
                      .IN8(na1873_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x138y38     80'h00_0018_00_0040_0C0F_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2290_1 ( .OUT(na2290_1), .IN1(na1843_1), .IN2(na1853_1), .IN3(na1863_1), .IN4(na1723_1), .IN5(na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x136y38     80'h00_0018_00_0040_0C0F_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2291_1 ( .OUT(na2291_1), .IN1(na2287_1), .IN2(na2288_1), .IN3(na2289_1), .IN4(na2290_1), .IN5(na2384_1), .IN6(1'b1), .IN7(na2385_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x154y40     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2292_1 ( .OUT(na2292_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1814_2), .IN6(na1734_2), .IN7(na1744_2),
                      .IN8(na1754_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x152y41     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2293_1 ( .OUT(na2293_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1794_2), .IN6(na1784_1), .IN7(na1774_2),
                      .IN8(na1764_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x153y36     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2294_1 ( .OUT(na2294_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1834_2), .IN6(na1824_2), .IN7(na1874_2),
                      .IN8(na1804_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x153y41     80'h00_0018_00_0040_0C0F_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2295_1 ( .OUT(na2295_1), .IN1(na1844_2), .IN2(na1854_1), .IN3(na1864_2), .IN4(na1724_2), .IN5(na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x148y40     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2296_1 ( .OUT(na2296_1), .IN1(~na2384_1), .IN2(1'b1), .IN3(~na2385_1), .IN4(1'b1), .IN5(na2295_1), .IN6(na2294_1), .IN7(na2293_1),
                      .IN8(na2292_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x140y43     80'h00_0018_00_0040_0C0F_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2297_1 ( .OUT(na2297_1), .IN1(na1745_1), .IN2(na1755_1), .IN3(na1815_1), .IN4(na1735_2), .IN5(na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x144y46     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2298_1 ( .OUT(na2298_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1775_1), .IN6(na1765_1), .IN7(na1795_1),
                      .IN8(na1785_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x143y43     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2299_1 ( .OUT(na2299_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1825_1), .IN6(na1835_1), .IN7(na1805_2),
                      .IN8(na1875_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x143y48     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2300_1 ( .OUT(na2300_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1725_1), .IN6(na1865_1), .IN7(na1855_1),
                      .IN8(na1845_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x138y50     80'h00_0018_00_0040_0C0F_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2301_1 ( .OUT(na2301_1), .IN1(na2299_1), .IN2(na2300_1), .IN3(na2297_1), .IN4(na2298_1), .IN5(na2384_1), .IN6(1'b1), .IN7(~na2385_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x152y46     80'h00_0018_00_0040_0C0F_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2302_1 ( .OUT(na2302_1), .IN1(na1816_2), .IN2(na1736_2), .IN3(na1746_2), .IN4(na1756_1), .IN5(na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x156y45     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2303_1 ( .OUT(na2303_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1766_2), .IN6(na1776_2), .IN7(na1786_2),
                      .IN8(na1796_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x153y48     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2304_1 ( .OUT(na2304_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1876_2), .IN6(na1806_2), .IN7(na1836_2),
                      .IN8(na1826_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x153y47     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2305_1 ( .OUT(na2305_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1856_2), .IN6(na1846_2), .IN7(na1726_2),
                      .IN8(na1866_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x154y50     80'h00_0018_00_0040_0C0F_5500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2306_1 ( .OUT(na2306_1), .IN1(na2305_1), .IN2(na2304_1), .IN3(na2303_1), .IN4(na2302_1), .IN5(~na2384_1), .IN6(1'b1), .IN7(~na2385_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x147y61     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2307_1 ( .OUT(na2307_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1737_1), .IN6(na1817_1), .IN7(na1757_1),
                      .IN8(na1747_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x153y62     80'h00_0018_00_0040_0C0F_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2308_1 ( .OUT(na2308_1), .IN1(na1767_1), .IN2(na1777_2), .IN3(na1787_1), .IN4(na1797_1), .IN5(na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x150y61     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2309_1 ( .OUT(na2309_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1837_1), .IN6(na1827_1), .IN7(na1877_1),
                      .IN8(na1807_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x152y62     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2310_1 ( .OUT(na2310_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1727_1), .IN6(na1867_1), .IN7(na1857_1),
                      .IN8(na1847_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x150y58     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2311_1 ( .OUT(na2311_1), .IN1(na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na2307_1), .IN6(na2308_1), .IN7(na2309_1),
                      .IN8(na2310_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x147y65     80'h00_0018_00_0040_0C0F_5500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2312_1 ( .OUT(na2312_1), .IN1(na1758_2), .IN2(na1748_2), .IN3(na1738_2), .IN4(na1818_2), .IN5(~na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x147y64     80'h00_0018_00_0040_0C0F_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2313_1 ( .OUT(na2313_1), .IN1(na1788_2), .IN2(na1798_1), .IN3(na1768_2), .IN4(na1778_2), .IN5(na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x152y65     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2314_1 ( .OUT(na2314_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1838_2), .IN6(na1828_2), .IN7(na1878_2),
                      .IN8(na1808_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x150y66     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2315_1 ( .OUT(na2315_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1858_2), .IN6(na1848_2), .IN7(na1728_1),
                      .IN8(na1868_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x148y64     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2316_1 ( .OUT(na2316_1), .IN1(na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na2312_1), .IN6(na2313_1), .IN7(na2314_1),
                      .IN8(na2315_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x151y65     80'h00_0018_00_0040_0C0F_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2317_1 ( .OUT(na2317_1), .IN1(na1819_2), .IN2(na1739_1), .IN3(na1749_2), .IN4(na1759_1), .IN5(na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x153y66     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2318_1 ( .OUT(na2318_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1769_1), .IN6(na1779_1), .IN7(na1789_1),
                      .IN8(na1799_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x154y69     80'h00_0018_00_0040_0C0F_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2319_1 ( .OUT(na2319_1), .IN1(na1809_1), .IN2(na1879_1), .IN3(na1829_1), .IN4(na1839_1), .IN5(na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x156y70     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2320_1 ( .OUT(na2320_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1859_1), .IN6(na1849_1), .IN7(na1729_1),
                      .IN8(na1869_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x154y66     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2321_1 ( .OUT(na2321_1), .IN1(na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na2317_1), .IN6(na2318_1), .IN7(na2319_1),
                      .IN8(na2320_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x153y78     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2322_1 ( .OUT(na2322_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1740_2), .IN6(na1820_2), .IN7(na1760_2),
                      .IN8(na1750_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x155y79     80'h00_0018_00_0040_0C0F_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2323_1 ( .OUT(na2323_1), .IN1(na1770_1), .IN2(na1780_2), .IN3(na1790_2), .IN4(na1800_2), .IN5(na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x156y78     80'h00_0018_00_0040_0C0F_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2324_1 ( .OUT(na2324_1), .IN1(na1880_2), .IN2(na1810_2), .IN3(na1840_1), .IN4(na1830_2), .IN5(~na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x154y81     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2325_1 ( .OUT(na2325_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1860_2), .IN6(na1850_2), .IN7(na1730_2),
                      .IN8(na1870_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x154y76     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2326_1 ( .OUT(na2326_1), .IN1(~na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na2323_1), .IN6(na2322_1), .IN7(na2325_1),
                      .IN8(na2324_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x141y77     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2327_1 ( .OUT(na2327_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na1761_1), .IN6(na1751_1), .IN7(na1741_1),
                      .IN8(na1821_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x139y76     80'h00_0018_00_0040_0C0F_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2328_1 ( .OUT(na2328_1), .IN1(na1771_1), .IN2(na1781_1), .IN3(na1791_2), .IN4(na1801_1), .IN5(na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x140y73     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2329_1 ( .OUT(na2329_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na1811_1), .IN6(na1881_1), .IN7(na1831_1),
                      .IN8(na1841_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x142y78     80'h00_0018_00_0040_0C0F_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2330_1 ( .OUT(na2330_1), .IN1(na1861_2), .IN2(na1851_1), .IN3(na1731_1), .IN4(na1871_1), .IN5(~na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x138y74     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2331_1 ( .OUT(na2331_1), .IN1(na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na2327_1), .IN6(na2328_1), .IN7(na2329_1),
                      .IN8(na2330_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x108y32     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2332_1 ( .OUT(na2332_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na482_1), .IN6(na472_2), .IN7(na462_2),
                      .IN8(na402_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x110y31     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2333_1 ( .OUT(na2333_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na492_2), .IN6(na512_2), .IN7(na532_1),
                      .IN8(na552_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x113y32     80'h00_0018_00_0040_0C0F_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2334_1 ( .OUT(na2334_1), .IN1(na572_2), .IN2(na442_2), .IN3(na582_2), .IN4(na562_1), .IN5(na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x111y31     80'h00_0018_00_0040_0C0F_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2335_1 ( .OUT(na2335_1), .IN1(na542_2), .IN2(na522_2), .IN3(na502_2), .IN4(na452_1), .IN5(na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x115y37     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2336_1 ( .OUT(na2336_1), .IN1(~na2384_1), .IN2(1'b1), .IN3(~na2385_1), .IN4(1'b1), .IN5(na2335_1), .IN6(na2334_1), .IN7(na2333_1),
                      .IN8(na2332_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x109y40     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2337_1 ( .OUT(na2337_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na403_1), .IN6(na463_2), .IN7(na473_1),
                      .IN8(na483_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x107y35     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2338_1 ( .OUT(na2338_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na493_2), .IN6(na513_1), .IN7(na533_1),
                      .IN8(na553_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x108y38     80'h00_0018_00_0040_0C0F_5500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2339_1 ( .OUT(na2339_1), .IN1(na563_1), .IN2(na583_1), .IN3(na443_1), .IN4(na573_2), .IN5(~na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x106y37     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2340_1 ( .OUT(na2340_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na543_2), .IN6(na523_1), .IN7(na503_1),
                      .IN8(na453_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x113y37     80'h00_0018_00_0040_0C0F_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2341_1 ( .OUT(na2341_1), .IN1(na2338_1), .IN2(na2337_1), .IN3(na2340_1), .IN4(na2339_1), .IN5(~na2384_1), .IN6(1'b1), .IN7(na2385_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x108y44     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2342_1 ( .OUT(na2342_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na404_2), .IN6(na464_2), .IN7(na474_1),
                      .IN8(na484_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x106y45     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2343_1 ( .OUT(na2343_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na554_1), .IN6(na534_2), .IN7(na514_2),
                      .IN8(na494_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x109y48     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2344_1 ( .OUT(na2344_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na574_2), .IN6(na444_1), .IN7(na584_1),
                      .IN8(na564_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x107y47     80'h00_0018_00_0040_0C0F_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2345_1 ( .OUT(na2345_1), .IN1(na544_2), .IN2(na524_2), .IN3(na504_1), .IN4(na454_2), .IN5(na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x105y46     80'h00_0018_00_0040_0C0F_5500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2346_1 ( .OUT(na2346_1), .IN1(na2345_1), .IN2(na2344_1), .IN3(na2343_1), .IN4(na2342_1), .IN5(~na2384_1), .IN6(1'b1), .IN7(~na2385_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x110y49     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2347_1 ( .OUT(na2347_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na405_2), .IN6(na465_1), .IN7(na475_1),
                      .IN8(na485_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x110y52     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2348_1 ( .OUT(na2348_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na535_1), .IN6(na555_1), .IN7(na495_1),
                      .IN8(na515_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x107y49     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2349_1 ( .OUT(na2349_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na575_1), .IN6(na445_1), .IN7(na585_1),
                      .IN8(na565_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x109y54     80'h00_0018_00_0040_0C0F_5500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2350_1 ( .OUT(na2350_1), .IN1(na455_2), .IN2(na505_1), .IN3(na525_1), .IN4(na545_1), .IN5(~na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x107y51     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2351_1 ( .OUT(na2351_1), .IN1(na2384_1), .IN2(1'b1), .IN3(~na2385_1), .IN4(1'b1), .IN5(na2349_1), .IN6(na2350_1), .IN7(na2347_1),
                      .IN8(na2348_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x109y53     80'h00_0018_00_0040_0C0F_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2352_1 ( .OUT(na2352_1), .IN1(na406_2), .IN2(na466_1), .IN3(na476_2), .IN4(na486_2), .IN5(na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x109y56     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2353_1 ( .OUT(na2353_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na536_2), .IN6(na556_2), .IN7(na496_1),
                      .IN8(na516_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x108y55     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2354_1 ( .OUT(na2354_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na586_2), .IN6(na566_2), .IN7(na576_1),
                      .IN8(na446_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x110y56     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2355_1 ( .OUT(na2355_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na526_1), .IN6(na546_2), .IN7(na456_2),
                      .IN8(na506_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x111y56     80'h00_0018_00_0040_0C0F_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2356_1 ( .OUT(na2356_1), .IN1(na2352_1), .IN2(na2353_1), .IN3(na2354_1), .IN4(na2355_1), .IN5(na2384_1), .IN6(1'b1), .IN7(na2385_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x109y61     80'h00_0018_00_0040_0C0F_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2357_1 ( .OUT(na2357_1), .IN1(na477_2), .IN2(na487_1), .IN3(na407_1), .IN4(na467_1), .IN5(na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x111y64     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2358_1 ( .OUT(na2358_1), .IN1(na2382_1), .IN2(1'b1), .IN3(~na2383_1), .IN4(1'b1), .IN5(na537_2), .IN6(na557_1), .IN7(na497_1),
                      .IN8(na517_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x112y63     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2359_1 ( .OUT(na2359_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na577_1), .IN6(na447_1), .IN7(na587_2),
                      .IN8(na567_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x112y66     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2360_1 ( .OUT(na2360_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na547_1), .IN6(na527_1), .IN7(na507_2),
                      .IN8(na457_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x113y62     80'h00_0018_00_0040_0C0F_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2361_1 ( .OUT(na2361_1), .IN1(na2357_1), .IN2(na2358_1), .IN3(na2359_1), .IN4(na2360_1), .IN5(na2384_1), .IN6(1'b1), .IN7(na2385_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x107y68     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2362_1 ( .OUT(na2362_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na468_2), .IN6(na408_1), .IN7(na488_1),
                      .IN8(na478_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x105y65     80'h00_0018_00_0040_0C0F_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2363_1 ( .OUT(na2363_1), .IN1(na538_2), .IN2(na558_2), .IN3(na498_2), .IN4(na518_1), .IN5(na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x110y70     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2364_1 ( .OUT(na2364_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na448_2), .IN6(na578_2), .IN7(na568_2),
                      .IN8(na588_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x110y67     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2365_1 ( .OUT(na2365_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na548_1), .IN6(na528_2), .IN7(na508_2),
                      .IN8(na458_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x113y66     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2366_1 ( .OUT(na2366_1), .IN1(~na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na2363_1), .IN6(na2362_1), .IN7(na2365_1),
                      .IN8(na2364_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x109y77     80'h00_0018_00_0040_0C0F_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2367_1 ( .OUT(na2367_1), .IN1(na409_1), .IN2(na469_1), .IN3(na479_1), .IN4(na489_1), .IN5(na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x107y76     80'h00_0018_00_0040_0C0F_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2368_1 ( .OUT(na2368_1), .IN1(na519_1), .IN2(na499_2), .IN3(na559_2), .IN4(na539_1), .IN5(~na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x110y81     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2369_1 ( .OUT(na2369_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na449_2), .IN6(na579_1), .IN7(na569_1),
                      .IN8(na589_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x110y80     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2370_1 ( .OUT(na2370_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na549_1), .IN6(na529_2), .IN7(na509_1),
                      .IN8(na459_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x109y76     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2371_1 ( .OUT(na2371_1), .IN1(na2384_1), .IN2(1'b1), .IN3(na2385_1), .IN4(1'b1), .IN5(na2367_1), .IN6(na2368_1), .IN7(na2369_1),
                      .IN8(na2370_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x110y71     80'h00_0018_00_0040_0C0F_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2372_1 ( .OUT(na2372_1), .IN1(na410_2), .IN2(na470_2), .IN3(na480_2), .IN4(na490_2), .IN5(na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x112y80     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2373_1 ( .OUT(na2373_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na520_2), .IN6(na500_2), .IN7(na560_2),
                      .IN8(na540_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x115y77     80'h00_0018_00_0040_0C0F_5500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2374_1 ( .OUT(na2374_1), .IN1(na570_1), .IN2(na590_2), .IN3(na450_2), .IN4(na580_2), .IN5(~na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x111y80     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2375_1 ( .OUT(na2375_1), .IN1(~na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na530_2), .IN6(na550_2), .IN7(na460_1),
                      .IN8(na510_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x114y73     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2376_1 ( .OUT(na2376_1), .IN1(na2384_1), .IN2(1'b1), .IN3(~na2385_1), .IN4(1'b1), .IN5(na2374_1), .IN6(na2375_1), .IN7(na2372_1),
                      .IN8(na2373_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x122y84     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2377_1 ( .OUT(na2377_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na411_2), .IN6(na471_2), .IN7(na481_1),
                      .IN8(na491_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x118y79     80'h00_0018_00_0040_0C0F_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2378_1 ( .OUT(na2378_1), .IN1(na541_1), .IN2(na561_1), .IN3(na501_1), .IN4(na521_2), .IN5(na2382_1), .IN6(1'b1), .IN7(~na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x121y78     80'h00_0018_00_0040_0C0F_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2379_1 ( .OUT(na2379_1), .IN1(na581_2), .IN2(na451_1), .IN3(na591_1), .IN4(na571_1), .IN5(na2382_1), .IN6(1'b1), .IN7(na2383_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x117y75     80'h00_0018_00_0040_0AF0_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2380_1 ( .OUT(na2380_1), .IN1(na2382_1), .IN2(1'b1), .IN3(na2383_1), .IN4(1'b1), .IN5(na551_2), .IN6(na531_1), .IN7(na511_1),
                      .IN8(na461_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x120y75     80'h00_0018_00_0040_0AF0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2381_1 ( .OUT(na2381_1), .IN1(~na2384_1), .IN2(1'b1), .IN3(~na2385_1), .IN4(1'b1), .IN5(na2380_1), .IN6(na2379_1), .IN7(na2378_1),
                      .IN8(na2377_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a2382 ( .Y(na2382_1), .I(addr[0]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a2383 ( .Y(na2383_1), .I(addr[1]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a2384 ( .Y(na2384_1), .I(addr[2]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a2385 ( .Y(na2385_1), .I(addr[3]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a2386 ( .Y(na2386_1), .I(addr[4]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a2387 ( .Y(na2387_1), .I(addr[5]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a2388 ( .Y(na2388_1), .I(addr[6]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a2389 ( .Y(na2389_1), .I(addr[7]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000090)) 
           _a2390 ( .Y(na2390_1), .I(clk) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a2391 ( .O(rdat[0]), .A(na2504_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a2392 ( .O(rdat[1]), .A(na2505_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a2393 ( .O(rdat[2]), .A(na2506_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a2394 ( .O(rdat[3]), .A(na2507_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a2395 ( .O(rdat[4]), .A(na2508_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a2396 ( .O(rdat[5]), .A(na2509_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a2397 ( .O(rdat[6]), .A(na2510_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a2398 ( .O(rdat[7]), .A(na2511_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a2399 ( .O(rdat[8]), .A(na2512_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a2400 ( .O(rdat[9]), .A(na2513_10) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a2401 ( .Y(na2401_1), .I(wdat[0]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a2402 ( .Y(na2402_1), .I(wdat[1]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a2403 ( .Y(na2403_1), .I(wdat[2]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a2404 ( .Y(na2404_1), .I(wdat[3]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a2405 ( .Y(na2405_1), .I(wdat[4]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a2406 ( .Y(na2406_1), .I(wdat[5]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a2407 ( .Y(na2407_1), .I(wdat[6]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a2408 ( .Y(na2408_1), .I(wdat[7]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a2409 ( .Y(na2409_1), .I(wdat[8]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a2410 ( .Y(na2410_1), .I(wdat[9]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a2411 ( .Y(na2411_1), .I(we) );
// C_AND///AND/      x130y45     80'h00_0078_00_0000_0C88_AACA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2412_1 ( .OUT(na2412_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na5_2), .IN6(1'b1), .IN7(na2036_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2412_4 ( .OUT(na2412_2), .IN1(na5_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1986_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x135y44     80'h00_0018_00_0000_0CEE_0700
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2413_1 ( .OUT(na2413_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2514_2), .IN6(~na2236_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
GLBOUT     #(.GLBOUT_CFG (64'h0000_0000_0000_0010)) 
           _a2414 ( .GLB0(na2414_1), .GLB1(_d3), .GLB2(_d4), .GLB3(_d5), .CLK_FB0(_d6), .CLK_FB1(_d7), .CLK_FB2(_d8), .CLK_FB3(_d9),
                    .CLK0_0(1'b0), .CLK0_90(1'b0), .CLK0_180(1'b0), .CLK0_270(1'b0), .CLK0_BYP(na2_1), .CLK1_0(1'b0), .CLK1_90(1'b0),
                    .CLK1_180(1'b0), .CLK1_270(1'b0), .CLK1_BYP(1'b0), .CLK2_0(1'b0), .CLK2_90(1'b0), .CLK2_180(1'b0), .CLK2_270(1'b0),
                    .CLK2_BYP(1'b0), .CLK3_0(1'b0), .CLK3_90(1'b0), .CLK3_180(1'b0), .CLK3_270(1'b0), .CLK3_BYP(1'b0), .USR_GLB0(1'b0),
                    .USR_GLB1(1'b0), .USR_GLB2(1'b0), .USR_GLB3(1'b0), .USR_FB0(1'b0), .USR_FB1(1'b0), .USR_FB2(1'b0), .USR_FB3(1'b0) );
// C_///OR/      x130y46     80'h00_0060_00_0000_0C0E_FF53
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a2415_4 ( .OUT(na2415_2), .IN1(1'b0), .IN2(~na2186_1), .IN3(~na7_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x132y44     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2416_1 ( .OUT(na2416_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na4_2), .IN7(1'b1), .IN8(na2086_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x122y61     80'h00_0060_00_0000_0C08_FF33
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2417_4 ( .OUT(na2417_2), .IN1(1'b1), .IN2(~na2386_1), .IN3(1'b1), .IN4(~na2388_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x144y44     80'h00_0078_00_0000_0C88_F8CA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2422_1 ( .OUT(na2422_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na13_2), .IN6(na1891_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2422_4 ( .OUT(na2422_2), .IN1(na13_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1941_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x131y48     80'h00_0018_00_0000_0CEE_0700
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2423_1 ( .OUT(na2423_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na5_1), .IN6(~na1991_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x131y47     80'h00_0060_00_0000_0C0E_FF35
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a2425_4 ( .OUT(na2425_2), .IN1(~na5_2), .IN2(1'b0), .IN3(1'b0), .IN4(~na2041_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x125y45     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2426_1 ( .OUT(na2426_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2517_2), .IN7(na2191_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x128y47     80'h00_0078_00_0000_0C88_F8AA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2431_1 ( .OUT(na2431_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na5_2), .IN6(na2046_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2431_4 ( .OUT(na2431_2), .IN1(na5_1), .IN2(1'b1), .IN3(na1996_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x129y50     80'h00_0060_00_0000_0C0E_FF33
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a2432_4 ( .OUT(na2432_2), .IN1(1'b0), .IN2(~na4_1), .IN3(1'b0), .IN4(~na2246_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x121y49     80'h00_0018_00_0000_0CEE_5300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2434_1 ( .OUT(na2434_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na2196_1), .IN7(~na7_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x131y43     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2435_4 ( .OUT(na2435_2), .IN1(na2096_1), .IN2(na4_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x136y54     80'h00_0078_00_0000_0C88_CAF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2440_1 ( .OUT(na2440_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na13_2), .IN6(1'b1), .IN7(1'b1), .IN8(na1901_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2440_4 ( .OUT(na2440_2), .IN1(na13_1), .IN2(na1951_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x126y49     80'h00_0018_00_0000_0CEE_3500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2441_1 ( .OUT(na2441_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na5_1), .IN6(1'b0), .IN7(1'b0), .IN8(~na2001_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x125y50     80'h00_0060_00_0000_0C0E_FF07
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a2443_4 ( .OUT(na2443_2), .IN1(~na2051_1), .IN2(~na2516_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x124y49     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2444_1 ( .OUT(na2444_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2201_1), .IN6(1'b1), .IN7(na7_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x122y52     80'h00_0078_00_0000_0C88_F8CA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2449_1 ( .OUT(na2449_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na5_2), .IN6(na2056_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2449_4 ( .OUT(na2449_2), .IN1(na5_1), .IN2(1'b1), .IN3(1'b1), .IN4(na2006_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x132y57     80'h00_0060_00_0000_0C0E_FF07
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a2450_4 ( .OUT(na2450_2), .IN1(~na2256_1), .IN2(~na4_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x125y53     80'h00_0018_00_0000_0CEE_7000
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2452_1 ( .OUT(na2452_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na7_1), .IN8(~na2206_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x128y52     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2453_4 ( .OUT(na2453_2), .IN1(na2106_1), .IN2(na4_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x124y55     80'h00_0078_00_0000_0C88_F8AA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2458_1 ( .OUT(na2458_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2111_1), .IN6(na4_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2458_4 ( .OUT(na2458_2), .IN1(na5_1), .IN2(1'b1), .IN3(na2011_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x137y58     80'h00_0018_00_0000_0CEE_5300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2459_1 ( .OUT(na2459_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na4_1), .IN7(~na2261_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x125y55     80'h00_0060_00_0000_0C0E_FF55
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a2461_4 ( .OUT(na2461_2), .IN1(~na5_2), .IN2(1'b0), .IN3(~na2061_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x125y59     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2462_1 ( .OUT(na2462_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na7_1), .IN8(na2211_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x129y64     80'h00_0078_00_0000_0C88_ACF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2467_1 ( .OUT(na2467_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na4_2), .IN7(na2116_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2467_4 ( .OUT(na2467_2), .IN1(na5_1), .IN2(na2016_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x127y61     80'h00_0060_00_0000_0C0E_FF33
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a2468_4 ( .OUT(na2468_2), .IN1(1'b0), .IN2(~na4_1), .IN3(1'b0), .IN4(~na2266_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x126y63     80'h00_0018_00_0000_0CEE_3500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2470_1 ( .OUT(na2470_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na5_2), .IN6(1'b0), .IN7(1'b0), .IN8(~na2066_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x122y63     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2471_4 ( .OUT(na2471_2), .IN1(1'b1), .IN2(1'b1), .IN3(na7_1), .IN4(na2216_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x124y63     80'h00_0078_00_0000_0C88_ACF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2476_1 ( .OUT(na2476_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na4_2), .IN7(na2121_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2476_4 ( .OUT(na2476_2), .IN1(na5_1), .IN2(na2021_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x136y64     80'h00_0018_00_0000_0CEE_0700
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2477_1 ( .OUT(na2477_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2271_1), .IN6(~na4_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x125y64     80'h00_0060_00_0000_0C0E_FF07
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a2479_4 ( .OUT(na2479_2), .IN1(~na2071_1), .IN2(~na2516_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x125y64     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2480_1 ( .OUT(na2480_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2221_1), .IN6(1'b1), .IN7(na7_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x126y66     80'h00_0078_00_0000_0C88_CACA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2485_1 ( .OUT(na2485_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na5_2), .IN6(1'b1), .IN7(1'b1), .IN8(na2076_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2485_4 ( .OUT(na2485_2), .IN1(na5_1), .IN2(1'b1), .IN3(1'b1), .IN4(na2026_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x140y69     80'h00_0060_00_0000_0C0E_FF07
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a2486_4 ( .OUT(na2486_2), .IN1(~na2515_2), .IN2(~na2276_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x127y68     80'h00_0018_00_0000_0CEE_5500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2488_1 ( .OUT(na2488_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2226_1), .IN6(1'b0), .IN7(~na7_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x140y65     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2489_4 ( .OUT(na2489_2), .IN1(1'b1), .IN2(na4_2), .IN3(1'b1), .IN4(na2126_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x135y68     80'h00_0078_00_0000_0C88_CAF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2494_1 ( .OUT(na2494_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na13_2), .IN6(1'b1), .IN7(1'b1), .IN8(na1931_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2494_4 ( .OUT(na2494_2), .IN1(na13_1), .IN2(na1981_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x130y65     80'h00_0018_00_0000_0CEE_5500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2495_1 ( .OUT(na2495_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na5_1), .IN6(1'b0), .IN7(~na2031_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x134y70     80'h00_0060_00_0000_0C0E_FF53
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a2497_4 ( .OUT(na2497_2), .IN1(1'b0), .IN2(~na2231_1), .IN3(~na7_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x134y66     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2498_1 ( .OUT(na2498_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na4_2), .IN7(na2131_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_Route1////      x130y58     80'h00_0018_00_0050_0C66_0000
C_Route1   #(.CPE_CFG (9'b0_0001_0000)) 
           _a2503_1 ( .OUT(na2503_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na279_4), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x160y27     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2504_4 ( .OUT(na2504_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a2504_6 ( .RAM_O2(na2504_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na2504_2), .COMP_OUT(1'b0) );
// C_///AND/      x160y31     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2505_4 ( .OUT(na2505_2), .IN1(na18_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a2505_6 ( .RAM_O2(na2505_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na2505_2), .COMP_OUT(1'b0) );
// C_///AND/      x160y35     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2506_4 ( .OUT(na2506_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na25_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a2506_6 ( .RAM_O2(na2506_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na2506_2), .COMP_OUT(1'b0) );
// C_///AND/      x160y39     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2507_4 ( .OUT(na2507_2), .IN1(1'b1), .IN2(1'b1), .IN3(na32_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a2507_6 ( .RAM_O2(na2507_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na2507_2), .COMP_OUT(1'b0) );
// C_///AND/      x160y43     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2508_4 ( .OUT(na2508_2), .IN1(1'b1), .IN2(1'b1), .IN3(na39_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a2508_6 ( .RAM_O2(na2508_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na2508_2), .COMP_OUT(1'b0) );
// C_///AND/      x160y47     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2509_4 ( .OUT(na2509_2), .IN1(na46_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a2509_6 ( .RAM_O2(na2509_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na2509_2), .COMP_OUT(1'b0) );
// C_///AND/      x160y51     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2510_4 ( .OUT(na2510_2), .IN1(na53_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a2510_6 ( .RAM_O2(na2510_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na2510_2), .COMP_OUT(1'b0) );
// C_///AND/      x160y55     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2511_4 ( .OUT(na2511_2), .IN1(1'b1), .IN2(na60_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a2511_6 ( .RAM_O2(na2511_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na2511_2), .COMP_OUT(1'b0) );
// C_///AND/      x160y59     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2512_4 ( .OUT(na2512_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na67_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a2512_6 ( .RAM_O2(na2512_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na2512_2), .COMP_OUT(1'b0) );
// C_///AND/      x160y69     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2513_4 ( .OUT(na2513_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na74_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a2513_6 ( .RAM_O2(na2513_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na2513_2), .COMP_OUT(1'b0) );
// C_////Bridge      x137y43     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2514_5 ( .OUT(na2514_2), .IN1(1'b0), .IN2(na4_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x141y69     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2515_5 ( .OUT(na2515_2), .IN1(1'b0), .IN2(na4_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x127y56     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2516_5 ( .OUT(na2516_2), .IN1(na5_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x127y46     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2517_5 ( .OUT(na2517_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na7_1), .IN8(1'b0) );
// C_////Bridge      x124y66     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2518_5 ( .OUT(na2518_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na10_1), .IN8(1'b0) );
// C_////Bridge      x121y59     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2519_5 ( .OUT(na2519_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na277_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x137y58     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2520_5 ( .OUT(na2520_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na277_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x137y56     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2521_5 ( .OUT(na2521_2), .IN1(1'b0), .IN2(1'b0), .IN3(na279_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x129y60     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2522_5 ( .OUT(na2522_2), .IN1(1'b0), .IN2(1'b0), .IN3(na279_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x133y51     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2523_5 ( .OUT(na2523_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na2449_1) );
// C_////Bridge      x134y57     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2524_5 ( .OUT(na2524_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na2503_1) );
endmodule
